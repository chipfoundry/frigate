VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2720.000 BY 2300.000 ;
  PIN gpio3_in[0]
    PORT
      LAYER met2 ;
        RECT 2657.050 2296.000 2657.330 2302.000 ;
    END
  END gpio3_in[0]
  PIN gpio3_in[1]
    PORT
      LAYER met2 ;
        RECT 2629.450 2296.000 2629.730 2302.000 ;
    END
  END gpio3_in[1]
  PIN gpio3_in[2]
    PORT
      LAYER met2 ;
        RECT 2601.850 2296.000 2602.130 2302.000 ;
    END
  END gpio3_in[2]
  PIN gpio3_in[3]
    PORT
      LAYER met2 ;
        RECT 2574.250 2296.000 2574.530 2302.000 ;
    END
  END gpio3_in[3]
  PIN gpio3_in[4]
    PORT
      LAYER met2 ;
        RECT 2546.650 2296.000 2546.930 2302.000 ;
    END
  END gpio3_in[4]
  PIN gpio3_in[5]
    PORT
      LAYER met2 ;
        RECT 2519.050 2296.000 2519.330 2302.000 ;
    END
  END gpio3_in[5]
  PIN gpio3_in[6]
    PORT
      LAYER met2 ;
        RECT 2491.450 2296.000 2491.730 2302.000 ;
    END
  END gpio3_in[6]
  PIN gpio3_in[7]
    PORT
      LAYER met2 ;
        RECT 2463.850 2296.000 2464.130 2302.000 ;
    END
  END gpio3_in[7]
  PIN gpio3_oeb[0]
    PORT
      LAYER met2 ;
        RECT 2638.650 2296.000 2638.930 2302.000 ;
    END
  END gpio3_oeb[0]
  PIN gpio3_oeb[1]
    PORT
      LAYER met2 ;
        RECT 2611.050 2296.000 2611.330 2302.000 ;
    END
  END gpio3_oeb[1]
  PIN gpio3_oeb[2]
    PORT
      LAYER met2 ;
        RECT 2583.450 2296.000 2583.730 2302.000 ;
    END
  END gpio3_oeb[2]
  PIN gpio3_oeb[3]
    PORT
      LAYER met2 ;
        RECT 2555.850 2296.000 2556.130 2302.000 ;
    END
  END gpio3_oeb[3]
  PIN gpio3_oeb[4]
    PORT
      LAYER met2 ;
        RECT 2528.250 2296.000 2528.530 2302.000 ;
    END
  END gpio3_oeb[4]
  PIN gpio3_oeb[5]
    PORT
      LAYER met2 ;
        RECT 2500.650 2296.000 2500.930 2302.000 ;
    END
  END gpio3_oeb[5]
  PIN gpio3_oeb[6]
    PORT
      LAYER met2 ;
        RECT 2473.050 2296.000 2473.330 2302.000 ;
    END
  END gpio3_oeb[6]
  PIN gpio3_oeb[7]
    PORT
      LAYER met2 ;
        RECT 2445.450 2296.000 2445.730 2302.000 ;
    END
  END gpio3_oeb[7]
  PIN gpio3_out[0]
    PORT
      LAYER met2 ;
        RECT 2647.850 2296.000 2648.130 2302.000 ;
    END
  END gpio3_out[0]
  PIN gpio3_out[1]
    PORT
      LAYER met2 ;
        RECT 2620.250 2296.000 2620.530 2302.000 ;
    END
  END gpio3_out[1]
  PIN gpio3_out[2]
    PORT
      LAYER met2 ;
        RECT 2592.650 2296.000 2592.930 2302.000 ;
    END
  END gpio3_out[2]
  PIN gpio3_out[3]
    PORT
      LAYER met2 ;
        RECT 2565.050 2296.000 2565.330 2302.000 ;
    END
  END gpio3_out[3]
  PIN gpio3_out[4]
    PORT
      LAYER met2 ;
        RECT 2537.450 2296.000 2537.730 2302.000 ;
    END
  END gpio3_out[4]
  PIN gpio3_out[5]
    PORT
      LAYER met2 ;
        RECT 2509.850 2296.000 2510.130 2302.000 ;
    END
  END gpio3_out[5]
  PIN gpio3_out[6]
    PORT
      LAYER met2 ;
        RECT 2482.250 2296.000 2482.530 2302.000 ;
    END
  END gpio3_out[6]
  PIN gpio3_out[7]
    PORT
      LAYER met2 ;
        RECT 2454.650 2296.000 2454.930 2302.000 ;
    END
  END gpio3_out[7]
  PIN gpio4_in[0]
    PORT
      LAYER met2 ;
        RECT 274.250 2296.000 274.530 2302.000 ;
    END
  END gpio4_in[0]
  PIN gpio4_in[1]
    PORT
      LAYER met2 ;
        RECT 246.650 2296.000 246.930 2302.000 ;
    END
  END gpio4_in[1]
  PIN gpio4_in[2]
    PORT
      LAYER met2 ;
        RECT 219.050 2296.000 219.330 2302.000 ;
    END
  END gpio4_in[2]
  PIN gpio4_in[3]
    PORT
      LAYER met2 ;
        RECT 191.450 2296.000 191.730 2302.000 ;
    END
  END gpio4_in[3]
  PIN gpio4_in[4]
    PORT
      LAYER met2 ;
        RECT 163.850 2296.000 164.130 2302.000 ;
    END
  END gpio4_in[4]
  PIN gpio4_in[5]
    PORT
      LAYER met2 ;
        RECT 136.250 2296.000 136.530 2302.000 ;
    END
  END gpio4_in[5]
  PIN gpio4_in[6]
    PORT
      LAYER met2 ;
        RECT 108.650 2296.000 108.930 2302.000 ;
    END
  END gpio4_in[6]
  PIN gpio4_in[7]
    PORT
      LAYER met2 ;
        RECT 81.050 2296.000 81.330 2302.000 ;
    END
  END gpio4_in[7]
  PIN gpio4_oeb[0]
    PORT
      LAYER met2 ;
        RECT 255.850 2296.000 256.130 2302.000 ;
    END
  END gpio4_oeb[0]
  PIN gpio4_oeb[1]
    PORT
      LAYER met2 ;
        RECT 228.250 2296.000 228.530 2302.000 ;
    END
  END gpio4_oeb[1]
  PIN gpio4_oeb[2]
    PORT
      LAYER met2 ;
        RECT 200.650 2296.000 200.930 2302.000 ;
    END
  END gpio4_oeb[2]
  PIN gpio4_oeb[3]
    PORT
      LAYER met2 ;
        RECT 173.050 2296.000 173.330 2302.000 ;
    END
  END gpio4_oeb[3]
  PIN gpio4_oeb[4]
    PORT
      LAYER met2 ;
        RECT 145.450 2296.000 145.730 2302.000 ;
    END
  END gpio4_oeb[4]
  PIN gpio4_oeb[5]
    PORT
      LAYER met2 ;
        RECT 117.850 2296.000 118.130 2302.000 ;
    END
  END gpio4_oeb[5]
  PIN gpio4_oeb[6]
    PORT
      LAYER met2 ;
        RECT 90.250 2296.000 90.530 2302.000 ;
    END
  END gpio4_oeb[6]
  PIN gpio4_oeb[7]
    PORT
      LAYER met2 ;
        RECT 62.650 2296.000 62.930 2302.000 ;
    END
  END gpio4_oeb[7]
  PIN gpio4_out[0]
    PORT
      LAYER met2 ;
        RECT 265.050 2296.000 265.330 2302.000 ;
    END
  END gpio4_out[0]
  PIN gpio4_out[1]
    PORT
      LAYER met2 ;
        RECT 237.450 2296.000 237.730 2302.000 ;
    END
  END gpio4_out[1]
  PIN gpio4_out[2]
    PORT
      LAYER met2 ;
        RECT 209.850 2296.000 210.130 2302.000 ;
    END
  END gpio4_out[2]
  PIN gpio4_out[3]
    PORT
      LAYER met2 ;
        RECT 182.250 2296.000 182.530 2302.000 ;
    END
  END gpio4_out[3]
  PIN gpio4_out[4]
    PORT
      LAYER met2 ;
        RECT 154.650 2296.000 154.930 2302.000 ;
    END
  END gpio4_out[4]
  PIN gpio4_out[5]
    PORT
      LAYER met2 ;
        RECT 127.050 2296.000 127.330 2302.000 ;
    END
  END gpio4_out[5]
  PIN gpio4_out[6]
    PORT
      LAYER met2 ;
        RECT 99.450 2296.000 99.730 2302.000 ;
    END
  END gpio4_out[6]
  PIN gpio4_out[7]
    PORT
      LAYER met2 ;
        RECT 71.850 2296.000 72.130 2302.000 ;
    END
  END gpio4_out[7]
  PIN HWDATA[18]
    PORT
      LAYER met2 ;
        RECT 649.110 -2.000 649.390 4.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    PORT
      LAYER met2 ;
        RECT 656.930 -2.000 657.210 4.000 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    PORT
      LAYER met2 ;
        RECT 516.170 -2.000 516.450 4.000 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    PORT
      LAYER met2 ;
        RECT 664.750 -2.000 665.030 4.000 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    PORT
      LAYER met2 ;
        RECT 672.570 -2.000 672.850 4.000 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    PORT
      LAYER met2 ;
        RECT 680.390 -2.000 680.670 4.000 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    PORT
      LAYER met2 ;
        RECT 688.210 -2.000 688.490 4.000 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    PORT
      LAYER met2 ;
        RECT 696.030 -2.000 696.310 4.000 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    PORT
      LAYER met2 ;
        RECT 703.850 -2.000 704.130 4.000 ;
    END
  END HWDATA[25]
  PIN HWDATA[2]
    PORT
      LAYER met2 ;
        RECT 523.990 -2.000 524.270 4.000 ;
    END
  END HWDATA[2]
  PIN HWDATA[3]
    PORT
      LAYER met2 ;
        RECT 531.810 -2.000 532.090 4.000 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    PORT
      LAYER met2 ;
        RECT 539.630 -2.000 539.910 4.000 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    PORT
      LAYER met2 ;
        RECT 547.450 -2.000 547.730 4.000 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    PORT
      LAYER met2 ;
        RECT 555.270 -2.000 555.550 4.000 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    PORT
      LAYER met2 ;
        RECT 563.090 -2.000 563.370 4.000 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    PORT
      LAYER met2 ;
        RECT 570.910 -2.000 571.190 4.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    PORT
      LAYER met2 ;
        RECT 578.730 -2.000 579.010 4.000 ;
    END
  END HWDATA[9]
  PIN HADDR[0]
    PORT
      LAYER met2 ;
        RECT 258.110 -2.000 258.390 4.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    PORT
      LAYER met2 ;
        RECT 336.310 -2.000 336.590 4.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    PORT
      LAYER met2 ;
        RECT 344.130 -2.000 344.410 4.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    PORT
      LAYER met2 ;
        RECT 351.950 -2.000 352.230 4.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    PORT
      LAYER met2 ;
        RECT 359.770 -2.000 360.050 4.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    PORT
      LAYER met2 ;
        RECT 367.590 -2.000 367.870 4.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    PORT
      LAYER met2 ;
        RECT 375.410 -2.000 375.690 4.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    PORT
      LAYER met2 ;
        RECT 383.230 -2.000 383.510 4.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    PORT
      LAYER met2 ;
        RECT 391.050 -2.000 391.330 4.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    PORT
      LAYER met2 ;
        RECT 398.870 -2.000 399.150 4.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    PORT
      LAYER met2 ;
        RECT 406.690 -2.000 406.970 4.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    PORT
      LAYER met2 ;
        RECT 265.930 -2.000 266.210 4.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    PORT
      LAYER met2 ;
        RECT 414.510 -2.000 414.790 4.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    PORT
      LAYER met2 ;
        RECT 422.330 -2.000 422.610 4.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    PORT
      LAYER met2 ;
        RECT 430.150 -2.000 430.430 4.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    PORT
      LAYER met2 ;
        RECT 437.970 -2.000 438.250 4.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    PORT
      LAYER met2 ;
        RECT 445.790 -2.000 446.070 4.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    PORT
      LAYER met2 ;
        RECT 453.610 -2.000 453.890 4.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    PORT
      LAYER met2 ;
        RECT 461.430 -2.000 461.710 4.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    PORT
      LAYER met2 ;
        RECT 469.250 -2.000 469.530 4.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    PORT
      LAYER met2 ;
        RECT 477.070 -2.000 477.350 4.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    PORT
      LAYER met2 ;
        RECT 484.890 -2.000 485.170 4.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    PORT
      LAYER met2 ;
        RECT 273.750 -2.000 274.030 4.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    PORT
      LAYER met2 ;
        RECT 492.710 -2.000 492.990 4.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    PORT
      LAYER met2 ;
        RECT 500.530 -2.000 500.810 4.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    PORT
      LAYER met2 ;
        RECT 281.570 -2.000 281.850 4.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    PORT
      LAYER met2 ;
        RECT 289.390 -2.000 289.670 4.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    PORT
      LAYER met2 ;
        RECT 297.210 -2.000 297.490 4.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    PORT
      LAYER met2 ;
        RECT 305.030 -2.000 305.310 4.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    PORT
      LAYER met2 ;
        RECT 312.850 -2.000 313.130 4.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    PORT
      LAYER met2 ;
        RECT 320.670 -2.000 320.950 4.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    PORT
      LAYER met2 ;
        RECT 328.490 -2.000 328.770 4.000 ;
    END
  END HADDR[9]
  PIN HCLK
    PORT
      LAYER met2 ;
        RECT 234.650 -2.000 234.930 4.000 ;
    END
  END HCLK
  PIN HRESETn
    PORT
      LAYER met2 ;
        RECT 242.470 -2.000 242.750 4.000 ;
    END
  END HRESETn
  PIN HSEL
    PORT
      LAYER met2 ;
        RECT 250.290 -2.000 250.570 4.000 ;
    END
  END HSEL
  PIN HWDATA[0]
    PORT
      LAYER met2 ;
        RECT 508.350 -2.000 508.630 4.000 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    PORT
      LAYER met2 ;
        RECT 586.550 -2.000 586.830 4.000 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    PORT
      LAYER met2 ;
        RECT 594.370 -2.000 594.650 4.000 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    PORT
      LAYER met2 ;
        RECT 602.190 -2.000 602.470 4.000 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    PORT
      LAYER met2 ;
        RECT 610.010 -2.000 610.290 4.000 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    PORT
      LAYER met2 ;
        RECT 617.830 -2.000 618.110 4.000 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    PORT
      LAYER met2 ;
        RECT 625.650 -2.000 625.930 4.000 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    PORT
      LAYER met2 ;
        RECT 633.470 -2.000 633.750 4.000 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    PORT
      LAYER met2 ;
        RECT 641.290 -2.000 641.570 4.000 ;
    END
  END HWDATA[17]
  PIN HRDATA[4]
    PORT
      LAYER met2 ;
        RECT 844.610 -2.000 844.890 4.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    PORT
      LAYER met2 ;
        RECT 852.430 -2.000 852.710 4.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    PORT
      LAYER met2 ;
        RECT 860.250 -2.000 860.530 4.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    PORT
      LAYER met2 ;
        RECT 868.070 -2.000 868.350 4.000 ;
    END
  END HRDATA[7]
  PIN HREADY
    PORT
      LAYER met2 ;
        RECT 758.590 -2.000 758.870 4.000 ;
    END
  END HREADY
  PIN HWDATA[27]
    PORT
      LAYER met2 ;
        RECT 719.490 -2.000 719.770 4.000 ;
    END
  END HWDATA[27]
  PIN HWRITE
    PORT
      LAYER met2 ;
        RECT 766.410 -2.000 766.690 4.000 ;
    END
  END HWRITE
  PIN HSIZE[0]
    PORT
      LAYER met2 ;
        RECT 789.870 -2.000 790.150 4.000 ;
    END
  END HSIZE[0]
  PIN HSIZE[1]
    PORT
      LAYER met2 ;
        RECT 797.690 -2.000 797.970 4.000 ;
    END
  END HSIZE[1]
  PIN HSIZE[2]
    PORT
      LAYER met2 ;
        RECT 805.510 -2.000 805.790 4.000 ;
    END
  END HSIZE[2]
  PIN HTRANS[0]
    PORT
      LAYER met2 ;
        RECT 774.230 -2.000 774.510 4.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    PORT
      LAYER met2 ;
        RECT 782.050 -2.000 782.330 4.000 ;
    END
  END HTRANS[1]
  PIN HWDATA[28]
    PORT
      LAYER met2 ;
        RECT 727.310 -2.000 727.590 4.000 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    PORT
      LAYER met2 ;
        RECT 735.130 -2.000 735.410 4.000 ;
    END
  END HWDATA[29]
  PIN HWDATA[26]
    PORT
      LAYER met2 ;
        RECT 711.670 -2.000 711.950 4.000 ;
    END
  END HWDATA[26]
  PIN HWDATA[30]
    PORT
      LAYER met2 ;
        RECT 742.950 -2.000 743.230 4.000 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    PORT
      LAYER met2 ;
        RECT 750.770 -2.000 751.050 4.000 ;
    END
  END HWDATA[31]
  PIN HRDATA[0]
    PORT
      LAYER met2 ;
        RECT 813.330 -2.000 813.610 4.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[1]
    PORT
      LAYER met2 ;
        RECT 821.150 -2.000 821.430 4.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[2]
    PORT
      LAYER met2 ;
        RECT 828.970 -2.000 829.250 4.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[3]
    PORT
      LAYER met2 ;
        RECT 836.790 -2.000 837.070 4.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[12]
    PORT
      LAYER met2 ;
        RECT 907.170 -2.000 907.450 4.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    PORT
      LAYER met2 ;
        RECT 914.990 -2.000 915.270 4.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    PORT
      LAYER met2 ;
        RECT 922.810 -2.000 923.090 4.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    PORT
      LAYER met2 ;
        RECT 930.630 -2.000 930.910 4.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    PORT
      LAYER met2 ;
        RECT 938.450 -2.000 938.730 4.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[8]
    PORT
      LAYER met2 ;
        RECT 875.890 -2.000 876.170 4.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    PORT
      LAYER met2 ;
        RECT 883.710 -2.000 883.990 4.000 ;
    END
  END HRDATA[9]
  PIN HRDATA[17]
    PORT
      LAYER met2 ;
        RECT 946.270 -2.000 946.550 4.000 ;
    END
  END HRDATA[17]
  PIN HREADYOUT
    PORT
      LAYER met2 ;
        RECT 1063.570 -2.000 1063.850 4.000 ;
    END
  END HREADYOUT
  PIN HRDATA[18]
    PORT
      LAYER met2 ;
        RECT 954.090 -2.000 954.370 4.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    PORT
      LAYER met2 ;
        RECT 961.910 -2.000 962.190 4.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[10]
    PORT
      LAYER met2 ;
        RECT 891.530 -2.000 891.810 4.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[20]
    PORT
      LAYER met2 ;
        RECT 969.730 -2.000 970.010 4.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    PORT
      LAYER met2 ;
        RECT 977.550 -2.000 977.830 4.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    PORT
      LAYER met2 ;
        RECT 985.370 -2.000 985.650 4.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    PORT
      LAYER met2 ;
        RECT 993.190 -2.000 993.470 4.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    PORT
      LAYER met2 ;
        RECT 1001.010 -2.000 1001.290 4.000 ;
    END
  END HRDATA[24]
  PIN user_irq[0]
    PORT
      LAYER met2 ;
        RECT 1071.390 -2.000 1071.670 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[10]
    PORT
      LAYER met2 ;
        RECT 1149.590 -2.000 1149.870 4.000 ;
    END
  END user_irq[10]
  PIN user_irq[11]
    PORT
      LAYER met2 ;
        RECT 1157.410 -2.000 1157.690 4.000 ;
    END
  END user_irq[11]
  PIN user_irq[12]
    PORT
      LAYER met2 ;
        RECT 1165.230 -2.000 1165.510 4.000 ;
    END
  END user_irq[12]
  PIN user_irq[13]
    PORT
      LAYER met2 ;
        RECT 1173.050 -2.000 1173.330 4.000 ;
    END
  END user_irq[13]
  PIN user_irq[14]
    PORT
      LAYER met2 ;
        RECT 1180.870 -2.000 1181.150 4.000 ;
    END
  END user_irq[14]
  PIN user_irq[15]
    PORT
      LAYER met2 ;
        RECT 1188.690 -2.000 1188.970 4.000 ;
    END
  END user_irq[15]
  PIN user_irq[1]
    PORT
      LAYER met2 ;
        RECT 1079.210 -2.000 1079.490 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    PORT
      LAYER met2 ;
        RECT 1087.030 -2.000 1087.310 4.000 ;
    END
  END user_irq[2]
  PIN user_irq[3]
    PORT
      LAYER met2 ;
        RECT 1094.850 -2.000 1095.130 4.000 ;
    END
  END user_irq[3]
  PIN user_irq[4]
    PORT
      LAYER met2 ;
        RECT 1102.670 -2.000 1102.950 4.000 ;
    END
  END user_irq[4]
  PIN user_irq[5]
    PORT
      LAYER met2 ;
        RECT 1110.490 -2.000 1110.770 4.000 ;
    END
  END user_irq[5]
  PIN user_irq[6]
    PORT
      LAYER met2 ;
        RECT 1118.310 -2.000 1118.590 4.000 ;
    END
  END user_irq[6]
  PIN user_irq[7]
    PORT
      LAYER met2 ;
        RECT 1126.130 -2.000 1126.410 4.000 ;
    END
  END user_irq[7]
  PIN user_irq[8]
    PORT
      LAYER met2 ;
        RECT 1133.950 -2.000 1134.230 4.000 ;
    END
  END user_irq[8]
  PIN user_irq[9]
    PORT
      LAYER met2 ;
        RECT 1141.770 -2.000 1142.050 4.000 ;
    END
  END user_irq[9]
  PIN HRDATA[25]
    PORT
      LAYER met2 ;
        RECT 1008.830 -2.000 1009.110 4.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    PORT
      LAYER met2 ;
        RECT 1016.650 -2.000 1016.930 4.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    PORT
      LAYER met2 ;
        RECT 1024.470 -2.000 1024.750 4.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    PORT
      LAYER met2 ;
        RECT 1032.290 -2.000 1032.570 4.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    PORT
      LAYER met2 ;
        RECT 1040.110 -2.000 1040.390 4.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[11]
    PORT
      LAYER met2 ;
        RECT 899.350 -2.000 899.630 4.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[30]
    PORT
      LAYER met2 ;
        RECT 1047.930 -2.000 1048.210 4.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    PORT
      LAYER met2 ;
        RECT 1055.750 -2.000 1056.030 4.000 ;
    END
  END HRDATA[31]
  PIN sio_oeb[1]
    PORT
      LAYER met2 ;
        RECT 2485.070 -2.000 2485.350 4.000 ;
    END
  END sio_oeb[1]
  PIN sio_out[0]
    PORT
      LAYER met2 ;
        RECT 2453.790 -2.000 2454.070 4.000 ;
    END
  END sio_out[0]
  PIN sio_out[1]
    PORT
      LAYER met2 ;
        RECT 2477.250 -2.000 2477.530 4.000 ;
    END
  END sio_out[1]
  PIN sio_in[0]
    PORT
      LAYER met2 ;
        RECT 2445.970 -2.000 2446.250 4.000 ;
    END
  END sio_in[0]
  PIN sio_in[1]
    PORT
      LAYER met2 ;
        RECT 2469.430 -2.000 2469.710 4.000 ;
    END
  END sio_in[1]
  PIN sio_oeb[0]
    PORT
      LAYER met2 ;
        RECT 2461.610 -2.000 2461.890 4.000 ;
    END
  END sio_oeb[0]
  PIN vssa1
    PORT
      LAYER met4 ;
        RECT 2621.510 0.000 2645.410 3.190 ;
    END
    PORT
      LAYER met4 ;
        RECT 2671.405 0.000 2695.305 3.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 2716.780 1842.855 2720.000 1866.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 2716.780 1892.750 2720.000 1916.650 ;
    END
  END vssa1
  PIN vdda1
    PORT
      LAYER met4 ;
        RECT 2551.405 0.000 2575.305 3.190 ;
    END
    PORT
      LAYER met4 ;
        RECT 2501.510 0.000 2525.410 3.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 2716.780 1772.755 2720.000 1796.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 2716.780 1722.860 2720.000 1746.760 ;
    END
  END vdda1
  PIN vdda2
    PORT
      LAYER met4 ;
        RECT 194.590 0.000 218.490 3.190 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.695 0.000 168.595 3.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1736.645 3.220 1760.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1786.540 3.220 1810.440 ;
    END
  END vdda2
  PIN vssa2
    PORT
      LAYER met4 ;
        RECT 24.695 0.000 48.595 3.190 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.590 0.000 98.490 3.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1851.645 3.220 1875.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1901.540 3.220 1925.440 ;
    END
  END vssa2
  PIN voutref
    PORT
      LAYER met4 ;
        RECT 1669.965 2298.500 1670.605 2300.000 ;
    END
  END voutref
  PIN ibias100
    PORT
      LAYER met4 ;
        RECT 1695.565 2298.500 1696.205 2300.000 ;
    END
  END ibias100
  PIN ibias50
    PORT
      LAYER met4 ;
        RECT 1693.005 2298.500 1693.645 2300.000 ;
    END
  END ibias50
  PIN gpio3_1_analog
    PORT
      LAYER met4 ;
        RECT 1749.325 2298.500 1749.965 2300.000 ;
    END
  END gpio3_1_analog
  PIN gpio3_2_analog
    PORT
      LAYER met4 ;
        RECT 1746.765 2298.500 1747.405 2300.000 ;
    END
  END gpio3_2_analog
  PIN gpio3_3_analog
    PORT
      LAYER met4 ;
        RECT 1744.205 2298.500 1744.845 2300.000 ;
    END
  END gpio3_3_analog
  PIN gpio3_4_analog
    PORT
      LAYER met4 ;
        RECT 1741.645 2298.500 1742.285 2300.000 ;
    END
  END gpio3_4_analog
  PIN gpio3_5_analog
    PORT
      LAYER met4 ;
        RECT 1739.085 2298.500 1739.725 2300.000 ;
    END
  END gpio3_5_analog
  PIN gpio3_6_analog
    PORT
      LAYER met4 ;
        RECT 1736.525 2298.500 1737.165 2300.000 ;
    END
  END gpio3_6_analog
  PIN gpio3_7_analog
    PORT
      LAYER met4 ;
        RECT 1733.965 2298.500 1734.605 2300.000 ;
    END
  END gpio3_7_analog
  PIN gpio4_0_analog
    PORT
      LAYER met4 ;
        RECT 1731.405 2298.500 1732.045 2300.000 ;
    END
  END gpio4_0_analog
  PIN gpio4_1_analog
    PORT
      LAYER met4 ;
        RECT 1728.845 2298.500 1729.485 2300.000 ;
    END
  END gpio4_1_analog
  PIN gpio4_2_analog
    PORT
      LAYER met4 ;
        RECT 1726.285 2298.500 1726.925 2300.000 ;
    END
  END gpio4_2_analog
  PIN gpio4_3_analog
    PORT
      LAYER met4 ;
        RECT 1723.725 2298.500 1724.365 2300.000 ;
    END
  END gpio4_3_analog
  PIN gpio4_4_analog
    PORT
      LAYER met4 ;
        RECT 1721.165 2298.500 1721.805 2300.000 ;
    END
  END gpio4_4_analog
  PIN gpio4_5_analog
    PORT
      LAYER met4 ;
        RECT 1718.605 2298.500 1719.245 2300.000 ;
    END
  END gpio4_5_analog
  PIN gpio4_6_analog
    PORT
      LAYER met4 ;
        RECT 1716.045 2298.500 1716.685 2300.000 ;
    END
  END gpio4_6_analog
  PIN gpio4_7_analog
    PORT
      LAYER met4 ;
        RECT 1713.485 2298.500 1714.125 2300.000 ;
    END
  END gpio4_7_analog
  PIN ulpcomp_p
    PORT
      LAYER met4 ;
        RECT 1710.925 2298.500 1711.565 2300.000 ;
    END
  END ulpcomp_p
  PIN ulpcomp_n
    PORT
      LAYER met4 ;
        RECT 1708.365 2298.500 1709.005 2300.000 ;
    END
  END ulpcomp_n
  PIN comp_p
    PORT
      LAYER met4 ;
        RECT 1705.805 2298.500 1706.445 2300.000 ;
    END
  END comp_p
  PIN comp_n
    PORT
      LAYER met4 ;
        RECT 1703.245 2298.500 1703.885 2300.000 ;
    END
  END comp_n
  PIN adc1
    PORT
      LAYER met4 ;
        RECT 1700.685 2298.500 1701.325 2300.000 ;
    END
  END adc1
  PIN adc0
    PORT
      LAYER met4 ;
        RECT 1698.125 2298.500 1698.765 2300.000 ;
    END
  END adc0
  PIN vbgsc
    PORT
      LAYER met4 ;
        RECT 1690.445 2298.500 1691.085 2300.000 ;
    END
  END vbgsc
  PIN vbgtc
    PORT
      LAYER met4 ;
        RECT 1687.885 2298.500 1688.525 2300.000 ;
    END
  END vbgtc
  PIN dac1
    PORT
      LAYER met4 ;
        RECT 1685.325 2298.500 1685.965 2300.000 ;
    END
  END dac1
  PIN dac0
    PORT
      LAYER met4 ;
        RECT 1682.765 2298.500 1683.405 2300.000 ;
    END
  END dac0
  PIN tempsense
    PORT
      LAYER met4 ;
        RECT 1680.205 2298.500 1680.845 2300.000 ;
    END
  END tempsense
  PIN right_vref
    PORT
      LAYER met4 ;
        RECT 1677.645 2298.500 1678.285 2300.000 ;
    END
  END right_vref
  PIN left_vref
    PORT
      LAYER met4 ;
        RECT 1675.085 2298.500 1675.725 2300.000 ;
    END
  END left_vref
  PIN vinref
    PORT
      LAYER met4 ;
        RECT 1672.525 2298.500 1673.165 2300.000 ;
    END
  END vinref
  PIN gpio3_0_analog
    PORT
      LAYER met4 ;
        RECT 1751.885 2298.500 1752.525 2300.000 ;
    END
  END gpio3_0_analog
  PIN gpio1_out[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 1264.840 2722.000 1265.440 ;
    END
  END gpio1_out[5]
  PIN gpio1_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 1287.960 2722.000 1288.560 ;
    END
  END gpio1_oeb[5]
  PIN gpio1_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 1357.320 2722.000 1357.920 ;
    END
  END gpio1_oeb[6]
  PIN gpio1_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 1426.680 2722.000 1427.280 ;
    END
  END gpio1_oeb[7]
  PIN gpio1_in[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 1311.080 2722.000 1311.680 ;
    END
  END gpio1_in[6]
  PIN gpio1_out[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 1334.200 2722.000 1334.800 ;
    END
  END gpio1_out[6]
  PIN gpio1_out[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 1403.560 2722.000 1404.160 ;
    END
  END gpio1_out[7]
  PIN gpio2_in[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 1449.800 2722.000 1450.400 ;
    END
  END gpio2_in[0]
  PIN gpio2_in[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 1519.160 2722.000 1519.760 ;
    END
  END gpio2_in[1]
  PIN gpio2_in[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 1588.520 2722.000 1589.120 ;
    END
  END gpio2_in[2]
  PIN gpio2_in[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 1657.880 2722.000 1658.480 ;
    END
  END gpio2_in[3]
  PIN gpio2_in[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 2027.800 2722.000 2028.400 ;
    END
  END gpio2_in[4]
  PIN gpio2_in[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 2097.160 2722.000 2097.760 ;
    END
  END gpio2_in[5]
  PIN gpio2_in[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 2166.520 2722.000 2167.120 ;
    END
  END gpio2_in[6]
  PIN gpio2_in[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 2235.880 2722.000 2236.480 ;
    END
  END gpio2_in[7]
  PIN gpio2_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 1496.040 2722.000 1496.640 ;
    END
  END gpio2_oeb[0]
  PIN gpio2_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 1565.400 2722.000 1566.000 ;
    END
  END gpio2_oeb[1]
  PIN gpio2_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 1634.760 2722.000 1635.360 ;
    END
  END gpio2_oeb[2]
  PIN gpio2_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 1704.120 2722.000 1704.720 ;
    END
  END gpio2_oeb[3]
  PIN gpio2_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 2074.040 2722.000 2074.640 ;
    END
  END gpio2_oeb[4]
  PIN gpio2_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 2143.400 2722.000 2144.000 ;
    END
  END gpio2_oeb[5]
  PIN gpio2_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 2212.760 2722.000 2213.360 ;
    END
  END gpio2_oeb[6]
  PIN gpio2_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 2282.120 2722.000 2282.720 ;
    END
  END gpio2_oeb[7]
  PIN gpio2_out[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 1472.920 2722.000 1473.520 ;
    END
  END gpio2_out[0]
  PIN gpio2_out[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 1542.280 2722.000 1542.880 ;
    END
  END gpio2_out[1]
  PIN gpio2_out[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 1611.640 2722.000 1612.240 ;
    END
  END gpio2_out[2]
  PIN gpio2_out[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 1681.000 2722.000 1681.600 ;
    END
  END gpio2_out[3]
  PIN gpio2_out[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 2050.920 2722.000 2051.520 ;
    END
  END gpio2_out[4]
  PIN gpio2_out[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 2120.280 2722.000 2120.880 ;
    END
  END gpio2_out[5]
  PIN gpio2_out[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 2189.640 2722.000 2190.240 ;
    END
  END gpio2_out[6]
  PIN gpio2_out[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 2259.000 2722.000 2259.600 ;
    END
  END gpio2_out[7]
  PIN gpio1_in[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 1380.440 2722.000 1381.040 ;
    END
  END gpio1_in[7]
  PIN gpio1_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 1218.600 2722.000 1219.200 ;
    END
  END gpio1_oeb[4]
  PIN gpio1_out[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 1195.480 2722.000 1196.080 ;
    END
  END gpio1_out[4]
  PIN gpio1_in[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 1241.720 2722.000 1242.320 ;
    END
  END gpio1_in[5]
  PIN gpio5_in[7]
    PORT
      LAYER met3 ;
        RECT -2.000 1496.040 4.000 1496.640 ;
    END
  END gpio5_in[7]
  PIN gpio5_oeb[0]
    PORT
      LAYER met3 ;
        RECT -2.000 2237.880 4.000 2238.480 ;
    END
  END gpio5_oeb[0]
  PIN gpio5_oeb[1]
    PORT
      LAYER met3 ;
        RECT -2.000 2168.520 4.000 2169.120 ;
    END
  END gpio5_oeb[1]
  PIN gpio5_oeb[2]
    PORT
      LAYER met3 ;
        RECT -2.000 2099.160 4.000 2099.760 ;
    END
  END gpio5_oeb[2]
  PIN gpio5_oeb[3]
    PORT
      LAYER met3 ;
        RECT -2.000 2029.800 4.000 2030.400 ;
    END
  END gpio5_oeb[3]
  PIN gpio5_oeb[4]
    PORT
      LAYER met3 ;
        RECT -2.000 1657.880 4.000 1658.480 ;
    END
  END gpio5_oeb[4]
  PIN gpio5_oeb[5]
    PORT
      LAYER met3 ;
        RECT -2.000 1588.520 4.000 1589.120 ;
    END
  END gpio5_oeb[5]
  PIN gpio5_oeb[6]
    PORT
      LAYER met3 ;
        RECT -2.000 1519.160 4.000 1519.760 ;
    END
  END gpio5_oeb[6]
  PIN gpio5_oeb[7]
    PORT
      LAYER met3 ;
        RECT -2.000 1449.800 4.000 1450.400 ;
    END
  END gpio5_oeb[7]
  PIN gpio5_out[0]
    PORT
      LAYER met3 ;
        RECT -2.000 2261.000 4.000 2261.600 ;
    END
  END gpio5_out[0]
  PIN gpio5_out[1]
    PORT
      LAYER met3 ;
        RECT -2.000 2191.640 4.000 2192.240 ;
    END
  END gpio5_out[1]
  PIN gpio5_out[2]
    PORT
      LAYER met3 ;
        RECT -2.000 2122.280 4.000 2122.880 ;
    END
  END gpio5_out[2]
  PIN gpio5_out[3]
    PORT
      LAYER met3 ;
        RECT -2.000 2052.920 4.000 2053.520 ;
    END
  END gpio5_out[3]
  PIN gpio5_out[4]
    PORT
      LAYER met3 ;
        RECT -2.000 1681.000 4.000 1681.600 ;
    END
  END gpio5_out[4]
  PIN gpio5_out[5]
    PORT
      LAYER met3 ;
        RECT -2.000 1611.640 4.000 1612.240 ;
    END
  END gpio5_out[5]
  PIN gpio5_out[6]
    PORT
      LAYER met3 ;
        RECT -2.000 1542.280 4.000 1542.880 ;
    END
  END gpio5_out[6]
  PIN gpio5_out[7]
    PORT
      LAYER met3 ;
        RECT -2.000 1472.920 4.000 1473.520 ;
    END
  END gpio5_out[7]
  PIN gpio6_in[0]
    PORT
      LAYER met3 ;
        RECT -2.000 1426.680 4.000 1427.280 ;
    END
  END gpio6_in[0]
  PIN gpio6_in[1]
    PORT
      LAYER met3 ;
        RECT -2.000 1357.320 4.000 1357.920 ;
    END
  END gpio6_in[1]
  PIN gpio6_in[2]
    PORT
      LAYER met3 ;
        RECT -2.000 1287.960 4.000 1288.560 ;
    END
  END gpio6_in[2]
  PIN gpio6_oeb[0]
    PORT
      LAYER met3 ;
        RECT -2.000 1380.440 4.000 1381.040 ;
    END
  END gpio6_oeb[0]
  PIN gpio6_oeb[1]
    PORT
      LAYER met3 ;
        RECT -2.000 1311.080 4.000 1311.680 ;
    END
  END gpio6_oeb[1]
  PIN gpio6_out[0]
    PORT
      LAYER met3 ;
        RECT -2.000 1403.560 4.000 1404.160 ;
    END
  END gpio6_out[0]
  PIN gpio6_out[1]
    PORT
      LAYER met3 ;
        RECT -2.000 1334.200 4.000 1334.800 ;
    END
  END gpio6_out[1]
  PIN gpio5_in[0]
    PORT
      LAYER met3 ;
        RECT -2.000 2284.120 4.000 2284.720 ;
    END
  END gpio5_in[0]
  PIN gpio5_in[1]
    PORT
      LAYER met3 ;
        RECT -2.000 2214.760 4.000 2215.360 ;
    END
  END gpio5_in[1]
  PIN gpio5_in[2]
    PORT
      LAYER met3 ;
        RECT -2.000 2145.400 4.000 2146.000 ;
    END
  END gpio5_in[2]
  PIN gpio5_in[3]
    PORT
      LAYER met3 ;
        RECT -2.000 2076.040 4.000 2076.640 ;
    END
  END gpio5_in[3]
  PIN gpio5_in[4]
    PORT
      LAYER met3 ;
        RECT -2.000 1704.120 4.000 1704.720 ;
    END
  END gpio5_in[4]
  PIN gpio6_out[3]
    PORT
      LAYER met3 ;
        RECT -2.000 1195.480 4.000 1196.080 ;
    END
  END gpio6_out[3]
  PIN gpio6_in[3]
    PORT
      LAYER met3 ;
        RECT -2.000 1218.600 4.000 1219.200 ;
    END
  END gpio6_in[3]
  PIN gpio6_oeb[2]
    PORT
      LAYER met3 ;
        RECT -2.000 1241.720 4.000 1242.320 ;
    END
  END gpio6_oeb[2]
  PIN gpio6_out[2]
    PORT
      LAYER met3 ;
        RECT -2.000 1264.840 4.000 1265.440 ;
    END
  END gpio6_out[2]
  PIN gpio5_in[5]
    PORT
      LAYER met3 ;
        RECT -2.000 1634.760 4.000 1635.360 ;
    END
  END gpio5_in[5]
  PIN gpio5_in[6]
    PORT
      LAYER met3 ;
        RECT -2.000 1565.400 4.000 1566.000 ;
    END
  END gpio5_in[6]
  PIN gpio6_out[6]
    PORT
      LAYER met3 ;
        RECT -2.000 987.400 4.000 988.000 ;
    END
  END gpio6_out[6]
  PIN gpio6_out[7]
    PORT
      LAYER met3 ;
        RECT -2.000 918.040 4.000 918.640 ;
    END
  END gpio6_out[7]
  PIN gpio7_in[0]
    PORT
      LAYER met3 ;
        RECT -2.000 870.320 4.000 870.920 ;
    END
  END gpio7_in[0]
  PIN gpio7_in[1]
    PORT
      LAYER met3 ;
        RECT -2.000 800.960 4.000 801.560 ;
    END
  END gpio7_in[1]
  PIN gpio7_in[2]
    PORT
      LAYER met3 ;
        RECT -2.000 731.600 4.000 732.200 ;
    END
  END gpio7_in[2]
  PIN gpio7_in[3]
    PORT
      LAYER met3 ;
        RECT -2.000 571.240 4.000 571.840 ;
    END
  END gpio7_in[3]
  PIN gpio7_in[4]
    PORT
      LAYER met3 ;
        RECT -2.000 501.880 4.000 502.480 ;
    END
  END gpio7_in[4]
  PIN gpio7_in[5]
    PORT
      LAYER met3 ;
        RECT -2.000 432.520 4.000 433.120 ;
    END
  END gpio7_in[5]
  PIN gpio7_in[6]
    PORT
      LAYER met3 ;
        RECT -2.000 363.160 4.000 363.760 ;
    END
  END gpio7_in[6]
  PIN gpio7_in[7]
    PORT
      LAYER met3 ;
        RECT -2.000 293.800 4.000 294.400 ;
    END
  END gpio7_in[7]
  PIN gpio7_oeb[0]
    PORT
      LAYER met3 ;
        RECT -2.000 824.080 4.000 824.680 ;
    END
  END gpio7_oeb[0]
  PIN gpio7_oeb[1]
    PORT
      LAYER met3 ;
        RECT -2.000 754.720 4.000 755.320 ;
    END
  END gpio7_oeb[1]
  PIN gpio7_oeb[2]
    PORT
      LAYER met3 ;
        RECT -2.000 594.360 4.000 594.960 ;
    END
  END gpio7_oeb[2]
  PIN gpio7_oeb[3]
    PORT
      LAYER met3 ;
        RECT -2.000 525.000 4.000 525.600 ;
    END
  END gpio7_oeb[3]
  PIN gpio7_oeb[4]
    PORT
      LAYER met3 ;
        RECT -2.000 455.640 4.000 456.240 ;
    END
  END gpio7_oeb[4]
  PIN gpio7_oeb[5]
    PORT
      LAYER met3 ;
        RECT -2.000 386.280 4.000 386.880 ;
    END
  END gpio7_oeb[5]
  PIN gpio7_oeb[6]
    PORT
      LAYER met3 ;
        RECT -2.000 316.920 4.000 317.520 ;
    END
  END gpio7_oeb[6]
  PIN gpio7_oeb[7]
    PORT
      LAYER met3 ;
        RECT -2.000 247.560 4.000 248.160 ;
    END
  END gpio7_oeb[7]
  PIN gpio7_out[0]
    PORT
      LAYER met3 ;
        RECT -2.000 847.200 4.000 847.800 ;
    END
  END gpio7_out[0]
  PIN gpio7_out[1]
    PORT
      LAYER met3 ;
        RECT -2.000 777.840 4.000 778.440 ;
    END
  END gpio7_out[1]
  PIN gpio7_out[2]
    PORT
      LAYER met3 ;
        RECT -2.000 617.480 4.000 618.080 ;
    END
  END gpio7_out[2]
  PIN gpio7_out[3]
    PORT
      LAYER met3 ;
        RECT -2.000 548.120 4.000 548.720 ;
    END
  END gpio7_out[3]
  PIN gpio7_out[4]
    PORT
      LAYER met3 ;
        RECT -2.000 478.760 4.000 479.360 ;
    END
  END gpio7_out[4]
  PIN gpio7_out[5]
    PORT
      LAYER met3 ;
        RECT -2.000 409.400 4.000 410.000 ;
    END
  END gpio7_out[5]
  PIN gpio7_out[6]
    PORT
      LAYER met3 ;
        RECT -2.000 340.040 4.000 340.640 ;
    END
  END gpio7_out[6]
  PIN gpio7_out[7]
    PORT
      LAYER met3 ;
        RECT -2.000 270.680 4.000 271.280 ;
    END
  END gpio7_out[7]
  PIN gpio6_in[6]
    PORT
      LAYER met3 ;
        RECT -2.000 1010.520 4.000 1011.120 ;
    END
  END gpio6_in[6]
  PIN gpio6_in[4]
    PORT
      LAYER met3 ;
        RECT -2.000 1149.240 4.000 1149.840 ;
    END
  END gpio6_in[4]
  PIN gpio6_in[7]
    PORT
      LAYER met3 ;
        RECT -2.000 941.160 4.000 941.760 ;
    END
  END gpio6_in[7]
  PIN gpio6_oeb[3]
    PORT
      LAYER met3 ;
        RECT -2.000 1172.360 4.000 1172.960 ;
    END
  END gpio6_oeb[3]
  PIN gpio6_oeb[4]
    PORT
      LAYER met3 ;
        RECT -2.000 1103.000 4.000 1103.600 ;
    END
  END gpio6_oeb[4]
  PIN gpio6_oeb[5]
    PORT
      LAYER met3 ;
        RECT -2.000 1033.640 4.000 1034.240 ;
    END
  END gpio6_oeb[5]
  PIN gpio6_oeb[6]
    PORT
      LAYER met3 ;
        RECT -2.000 964.280 4.000 964.880 ;
    END
  END gpio6_oeb[6]
  PIN gpio6_oeb[7]
    PORT
      LAYER met3 ;
        RECT -2.000 894.920 4.000 895.520 ;
    END
  END gpio6_oeb[7]
  PIN gpio6_in[5]
    PORT
      LAYER met3 ;
        RECT -2.000 1079.880 4.000 1080.480 ;
    END
  END gpio6_in[5]
  PIN gpio6_out[4]
    PORT
      LAYER met3 ;
        RECT -2.000 1126.120 4.000 1126.720 ;
    END
  END gpio6_out[4]
  PIN gpio6_out[5]
    PORT
      LAYER met3 ;
        RECT -2.000 1056.760 4.000 1057.360 ;
    END
  END gpio6_out[5]
  PIN gpio1_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 1149.240 2722.000 1149.840 ;
    END
  END gpio1_oeb[3]
  PIN gpio1_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 941.160 2722.000 941.760 ;
    END
  END gpio1_oeb[0]
  PIN gpio0_in[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 235.810 2722.000 236.410 ;
    END
  END gpio0_in[2]
  PIN gpio0_in[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 305.170 2722.000 305.770 ;
    END
  END gpio0_in[3]
  PIN gpio0_in[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 374.530 2722.000 375.130 ;
    END
  END gpio0_in[4]
  PIN gpio1_out[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 918.040 2722.000 918.640 ;
    END
  END gpio1_out[0]
  PIN gpio1_out[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 987.400 2722.000 988.000 ;
    END
  END gpio1_out[1]
  PIN gpio1_out[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 1056.760 2722.000 1057.360 ;
    END
  END gpio1_out[2]
  PIN gpio1_out[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 1126.120 2722.000 1126.720 ;
    END
  END gpio1_out[3]
  PIN gpio1_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 1010.520 2722.000 1011.120 ;
    END
  END gpio1_oeb[1]
  PIN gpio0_in[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 443.890 2722.000 444.490 ;
    END
  END gpio0_in[5]
  PIN gpio0_in[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 513.250 2722.000 513.850 ;
    END
  END gpio0_in[6]
  PIN gpio0_in[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 582.610 2722.000 583.210 ;
    END
  END gpio0_in[7]
  PIN gpio0_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 143.330 2722.000 143.930 ;
    END
  END gpio0_oeb[0]
  PIN gpio0_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 212.690 2722.000 213.290 ;
    END
  END gpio0_oeb[1]
  PIN gpio0_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 282.050 2722.000 282.650 ;
    END
  END gpio0_oeb[2]
  PIN gpio0_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 351.410 2722.000 352.010 ;
    END
  END gpio0_oeb[3]
  PIN gpio0_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 420.770 2722.000 421.370 ;
    END
  END gpio0_oeb[4]
  PIN gpio0_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 490.130 2722.000 490.730 ;
    END
  END gpio0_oeb[5]
  PIN gpio0_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 559.490 2722.000 560.090 ;
    END
  END gpio0_oeb[6]
  PIN gpio0_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 628.850 2722.000 629.450 ;
    END
  END gpio0_oeb[7]
  PIN gpio0_out[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 120.210 2722.000 120.810 ;
    END
  END gpio0_out[0]
  PIN gpio0_out[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 189.570 2722.000 190.170 ;
    END
  END gpio0_out[1]
  PIN gpio0_out[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 258.930 2722.000 259.530 ;
    END
  END gpio0_out[2]
  PIN gpio0_out[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 328.290 2722.000 328.890 ;
    END
  END gpio0_out[3]
  PIN gpio0_out[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 397.650 2722.000 398.250 ;
    END
  END gpio0_out[4]
  PIN gpio0_out[5]
    PORT
      LAYER met3 ;
        RECT 2716.000 467.010 2722.000 467.610 ;
    END
  END gpio0_out[5]
  PIN gpio0_out[6]
    PORT
      LAYER met3 ;
        RECT 2716.000 536.370 2722.000 536.970 ;
    END
  END gpio0_out[6]
  PIN gpio0_out[7]
    PORT
      LAYER met3 ;
        RECT 2716.000 605.730 2722.000 606.330 ;
    END
  END gpio0_out[7]
  PIN gpio1_in[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 894.920 2722.000 895.520 ;
    END
  END gpio1_in[0]
  PIN gpio1_in[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 964.280 2722.000 964.880 ;
    END
  END gpio1_in[1]
  PIN gpio1_in[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 1033.640 2722.000 1034.240 ;
    END
  END gpio1_in[2]
  PIN gpio1_in[3]
    PORT
      LAYER met3 ;
        RECT 2716.000 1103.000 2722.000 1103.600 ;
    END
  END gpio1_in[3]
  PIN gpio1_in[4]
    PORT
      LAYER met3 ;
        RECT 2716.000 1172.360 2722.000 1172.960 ;
    END
  END gpio1_in[4]
  PIN gpio1_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2716.000 1079.880 2722.000 1080.480 ;
    END
  END gpio1_oeb[2]
  PIN gpio0_in[0]
    PORT
      LAYER met3 ;
        RECT 2716.000 97.090 2722.000 97.690 ;
    END
  END gpio0_in[0]
  PIN gpio0_in[1]
    PORT
      LAYER met3 ;
        RECT 2716.000 166.450 2722.000 167.050 ;
    END
  END gpio0_in[1]
  OBS
      LAYER met2 ;
        RECT 6.530 710.075 6.810 710.445 ;
        RECT 6.600 708.890 6.740 710.075 ;
        RECT 6.540 708.570 6.800 708.890 ;
        RECT 6.530 640.715 6.810 641.085 ;
        RECT 6.540 640.570 6.800 640.715 ;
  END
END user_project_wrapper
END LIBRARY

