VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO product_id_rom_8bit
  CLASS BLOCK ;
  FOREIGN product_id_rom_8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.020 BY 11.000 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 10.135 8.350 10.565 9.135 ;
        RECT 14.195 8.350 14.625 9.135 ;
        RECT 14.195 7.185 14.625 7.970 ;
        RECT 10.135 2.910 10.565 3.695 ;
        RECT 14.195 2.910 14.625 3.695 ;
      LAYER li1 ;
        RECT 0.085 8.995 0.605 9.535 ;
        RECT 1.465 9.015 2.675 9.535 ;
        RECT 4.225 9.015 6.805 9.535 ;
        RECT 10.665 9.015 11.875 9.535 ;
        RECT 0.085 8.245 1.295 8.995 ;
        RECT 1.465 8.245 4.055 9.015 ;
        RECT 4.225 8.245 9.570 9.015 ;
        RECT 10.205 8.245 10.495 8.970 ;
        RECT 10.665 8.245 13.255 9.015 ;
        RECT 15.415 8.995 15.935 9.535 ;
        RECT 14.265 8.245 14.555 8.970 ;
        RECT 14.725 8.245 15.935 8.995 ;
        RECT 0.000 8.075 13.800 8.245 ;
        RECT 14.180 8.075 16.020 8.245 ;
        RECT 0.085 7.325 1.295 8.075 ;
        RECT 0.085 6.785 0.605 7.325 ;
        RECT 1.465 7.305 4.055 8.075 ;
        RECT 4.225 7.305 9.570 8.075 ;
        RECT 9.745 7.305 12.335 8.075 ;
        RECT 12.505 7.325 13.715 8.075 ;
        RECT 14.265 7.350 14.555 8.075 ;
        RECT 14.725 7.325 15.935 8.075 ;
        RECT 1.465 6.785 2.675 7.305 ;
        RECT 4.225 6.785 6.805 7.305 ;
        RECT 9.745 6.785 10.955 7.305 ;
        RECT 13.195 6.785 13.715 7.325 ;
        RECT 15.415 6.785 15.935 7.325 ;
        RECT 0.085 3.555 0.605 4.095 ;
        RECT 15.415 3.555 15.935 4.095 ;
        RECT 0.085 2.805 1.295 3.555 ;
        RECT 2.615 2.805 2.955 3.465 ;
        RECT 3.995 2.805 4.335 3.465 ;
        RECT 5.375 2.805 5.715 3.465 ;
        RECT 6.755 2.805 7.095 3.465 ;
        RECT 8.135 2.805 8.475 3.465 ;
        RECT 9.515 2.805 9.855 3.465 ;
        RECT 10.205 2.805 10.495 3.530 ;
        RECT 11.815 2.805 12.155 3.465 ;
        RECT 13.195 2.805 13.535 3.465 ;
        RECT 14.265 2.805 14.555 3.530 ;
        RECT 14.725 2.805 15.935 3.555 ;
        RECT 0.000 2.635 13.800 2.805 ;
        RECT 14.180 2.635 16.020 2.805 ;
      LAYER met1 ;
        RECT 0.000 7.920 16.020 8.400 ;
        RECT 0.000 2.480 16.020 2.960 ;
      LAYER met2 ;
        RECT 1.130 7.920 2.350 8.400 ;
        RECT 8.130 7.920 9.350 8.400 ;
        RECT 1.290 2.960 1.830 7.920 ;
        RECT 1.130 2.480 2.350 2.960 ;
        RECT 8.130 2.480 9.350 2.960 ;
      LAYER met3 ;
        RECT 1.040 7.920 9.440 8.400 ;
        RECT 1.040 2.480 9.440 2.960 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 9.465 16.210 11.070 ;
        RECT -0.190 4.025 16.210 6.855 ;
      LAYER li1 ;
        RECT 0.000 10.795 13.800 10.965 ;
        RECT 14.180 10.795 16.020 10.965 ;
        RECT 0.085 9.705 1.295 10.795 ;
        RECT 1.465 9.705 4.055 10.795 ;
        RECT 4.225 9.705 9.570 10.795 ;
        RECT 0.775 9.165 1.295 9.705 ;
        RECT 2.845 9.185 4.055 9.705 ;
        RECT 6.975 9.185 9.570 9.705 ;
        RECT 10.205 9.630 10.495 10.795 ;
        RECT 10.665 9.705 13.255 10.795 ;
        RECT 12.045 9.185 13.255 9.705 ;
        RECT 14.265 9.630 14.555 10.795 ;
        RECT 14.725 9.705 15.935 10.795 ;
        RECT 14.725 9.165 15.245 9.705 ;
        RECT 0.775 6.615 1.295 7.155 ;
        RECT 2.845 6.615 4.055 7.135 ;
        RECT 6.975 6.615 9.570 7.135 ;
        RECT 11.125 6.615 12.335 7.135 ;
        RECT 0.085 5.525 1.295 6.615 ;
        RECT 1.465 5.525 4.055 6.615 ;
        RECT 4.225 5.525 9.570 6.615 ;
        RECT 9.745 5.525 12.335 6.615 ;
        RECT 12.505 6.615 13.025 7.155 ;
        RECT 12.505 5.525 13.715 6.615 ;
        RECT 14.265 5.525 14.555 6.690 ;
        RECT 14.725 6.615 15.245 7.155 ;
        RECT 14.725 5.525 15.935 6.615 ;
        RECT 0.000 5.355 13.800 5.525 ;
        RECT 14.180 5.355 16.020 5.525 ;
        RECT 0.085 4.265 1.295 5.355 ;
        RECT 2.115 4.630 2.445 5.355 ;
        RECT 3.495 4.630 3.825 5.355 ;
        RECT 4.875 4.630 5.205 5.355 ;
        RECT 6.255 4.630 6.585 5.355 ;
        RECT 7.635 4.630 7.965 5.355 ;
        RECT 9.015 4.630 9.345 5.355 ;
        RECT 0.775 3.725 1.295 4.265 ;
        RECT 10.205 4.190 10.495 5.355 ;
        RECT 11.315 4.630 11.645 5.355 ;
        RECT 12.695 4.630 13.025 5.355 ;
        RECT 14.265 4.190 14.555 5.355 ;
        RECT 14.725 4.265 15.935 5.355 ;
        RECT 14.725 3.725 15.245 4.265 ;
      LAYER met1 ;
        RECT 0.000 10.640 16.020 11.120 ;
        RECT 0.000 5.200 16.020 5.680 ;
      LAYER met2 ;
        RECT 4.630 10.640 5.850 11.120 ;
        RECT 11.630 10.640 12.850 11.120 ;
        RECT 4.990 5.680 5.530 10.640 ;
        RECT 4.630 5.200 5.850 5.680 ;
        RECT 11.630 5.200 12.850 5.680 ;
      LAYER met3 ;
        RECT 4.540 10.640 12.940 11.120 ;
        RECT 4.540 5.200 12.940 5.680 ;
    END
  END VPWR
  PIN gpio_defaults[0]
    PORT
      LAYER li1 ;
        RECT 2.615 3.635 3.135 5.185 ;
      LAYER met1 ;
        RECT 2.035 3.980 2.325 4.025 ;
        RECT 2.725 3.980 3.015 4.025 ;
        RECT 2.035 3.840 3.015 3.980 ;
        RECT 2.035 3.795 2.325 3.840 ;
        RECT 2.725 3.795 3.015 3.840 ;
        RECT 2.815 3.555 2.955 3.795 ;
        RECT 2.770 3.235 3.030 3.555 ;
      LAYER met2 ;
        RECT 2.740 3.465 3.060 3.525 ;
        RECT 2.610 3.265 3.060 3.465 ;
        RECT 2.610 2.370 2.750 3.265 ;
        RECT 2.455 2.225 2.750 2.370 ;
        RECT 2.455 2.000 2.595 2.225 ;
        RECT 2.390 0.000 2.670 2.000 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[1]
    PORT
      LAYER li1 ;
        RECT 3.995 3.635 4.515 5.185 ;
      LAYER met1 ;
        RECT 3.415 3.980 3.705 4.025 ;
        RECT 4.105 3.980 4.395 4.025 ;
        RECT 3.415 3.840 4.395 3.980 ;
        RECT 3.415 3.795 3.705 3.840 ;
        RECT 4.105 3.795 4.395 3.840 ;
        RECT 4.195 3.555 4.335 3.795 ;
        RECT 4.150 3.235 4.410 3.555 ;
      LAYER met2 ;
        RECT 4.120 3.465 4.440 3.525 ;
        RECT 3.840 3.325 4.440 3.465 ;
        RECT 3.840 2.000 3.980 3.325 ;
        RECT 4.120 3.265 4.440 3.325 ;
        RECT 3.770 0.000 4.050 2.000 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[2]
    PORT
      LAYER li1 ;
        RECT 5.375 3.635 5.895 5.185 ;
      LAYER met1 ;
        RECT 4.795 3.980 5.085 4.025 ;
        RECT 5.485 3.980 5.775 4.025 ;
        RECT 4.795 3.840 5.775 3.980 ;
        RECT 4.795 3.795 5.085 3.840 ;
        RECT 5.485 3.795 5.775 3.840 ;
        RECT 5.575 3.555 5.715 3.795 ;
        RECT 5.530 3.235 5.790 3.555 ;
      LAYER met2 ;
        RECT 5.500 3.465 5.820 3.525 ;
        RECT 5.220 3.325 5.820 3.465 ;
        RECT 5.220 2.000 5.360 3.325 ;
        RECT 5.500 3.265 5.820 3.325 ;
        RECT 5.150 0.000 5.430 2.000 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[3]
    PORT
      LAYER li1 ;
        RECT 6.755 3.635 7.275 5.185 ;
      LAYER met1 ;
        RECT 6.175 3.980 6.465 4.025 ;
        RECT 6.865 3.980 7.155 4.025 ;
        RECT 6.175 3.840 7.155 3.980 ;
        RECT 6.175 3.795 6.465 3.840 ;
        RECT 6.865 3.795 7.155 3.840 ;
        RECT 6.955 3.555 7.095 3.795 ;
        RECT 6.910 3.235 7.170 3.555 ;
      LAYER met2 ;
        RECT 6.880 3.465 7.200 3.525 ;
        RECT 6.600 3.325 7.200 3.465 ;
        RECT 6.600 2.000 6.740 3.325 ;
        RECT 6.880 3.265 7.200 3.325 ;
        RECT 6.530 0.000 6.810 2.000 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[4]
    PORT
      LAYER li1 ;
        RECT 8.135 3.635 8.655 5.185 ;
      LAYER met1 ;
        RECT 7.555 3.980 7.845 4.025 ;
        RECT 8.245 3.980 8.535 4.025 ;
        RECT 7.555 3.840 8.535 3.980 ;
        RECT 7.555 3.795 7.845 3.840 ;
        RECT 8.245 3.795 8.535 3.840 ;
        RECT 8.335 3.555 8.475 3.795 ;
        RECT 8.290 3.235 8.550 3.555 ;
      LAYER met2 ;
        RECT 8.260 3.465 8.580 3.525 ;
        RECT 7.780 3.325 8.580 3.465 ;
        RECT 7.780 2.325 7.920 3.325 ;
        RECT 8.260 3.265 8.580 3.325 ;
        RECT 7.780 2.185 8.120 2.325 ;
        RECT 7.980 2.000 8.120 2.185 ;
        RECT 7.910 0.000 8.190 2.000 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[5]
    PORT
      LAYER li1 ;
        RECT 9.515 3.635 10.035 5.185 ;
      LAYER met1 ;
        RECT 8.935 3.980 9.225 4.025 ;
        RECT 9.625 3.980 9.915 4.025 ;
        RECT 8.935 3.840 9.915 3.980 ;
        RECT 8.935 3.795 9.225 3.840 ;
        RECT 9.625 3.795 9.915 3.840 ;
        RECT 9.715 3.555 9.855 3.795 ;
        RECT 9.670 3.235 9.930 3.555 ;
      LAYER met2 ;
        RECT 9.640 3.265 9.960 3.525 ;
        RECT 9.725 2.415 9.865 3.265 ;
        RECT 9.725 2.265 9.960 2.415 ;
        RECT 9.820 2.000 9.960 2.265 ;
        RECT 9.750 0.000 10.030 2.000 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[6]
    PORT
      LAYER li1 ;
        RECT 11.815 3.635 12.335 5.185 ;
      LAYER met1 ;
        RECT 11.235 3.980 11.525 4.025 ;
        RECT 11.925 3.980 12.215 4.025 ;
        RECT 11.235 3.840 12.215 3.980 ;
        RECT 11.235 3.795 11.525 3.840 ;
        RECT 11.925 3.795 12.215 3.840 ;
        RECT 12.015 3.555 12.155 3.795 ;
        RECT 11.970 3.235 12.230 3.555 ;
      LAYER met2 ;
        RECT 11.940 3.465 12.260 3.525 ;
        RECT 11.660 3.325 12.260 3.465 ;
        RECT 11.660 2.000 11.800 3.325 ;
        RECT 11.940 3.265 12.260 3.325 ;
        RECT 11.590 0.000 11.870 2.000 ;
    END
  END gpio_defaults[6]
  PIN gpio_defaults[7]
    PORT
      LAYER li1 ;
        RECT 13.195 3.635 13.715 5.185 ;
      LAYER met1 ;
        RECT 12.615 3.980 12.905 4.025 ;
        RECT 13.305 3.980 13.595 4.025 ;
        RECT 12.615 3.840 13.595 3.980 ;
        RECT 12.615 3.795 12.905 3.840 ;
        RECT 13.305 3.795 13.595 3.840 ;
        RECT 13.395 3.555 13.535 3.795 ;
        RECT 13.350 3.235 13.610 3.555 ;
      LAYER met2 ;
        RECT 13.320 3.465 13.640 3.525 ;
        RECT 13.040 3.325 13.640 3.465 ;
        RECT 13.040 2.000 13.180 3.325 ;
        RECT 13.320 3.265 13.640 3.325 ;
        RECT 12.970 0.000 13.250 2.000 ;
    END
  END gpio_defaults[7]
  OBS
      LAYER pwell ;
        RECT 0.005 8.265 1.375 9.075 ;
        RECT 1.385 8.265 4.135 9.075 ;
        RECT 4.145 8.265 9.655 9.075 ;
        RECT 10.585 8.265 13.335 9.075 ;
        RECT 14.645 8.265 16.015 9.075 ;
        RECT 0.145 8.055 0.315 8.265 ;
        RECT 1.525 8.055 1.695 8.265 ;
        RECT 4.285 8.055 4.455 8.265 ;
        RECT 9.805 8.215 9.975 8.245 ;
        RECT 9.800 8.105 9.975 8.215 ;
        RECT 9.805 8.055 9.975 8.105 ;
        RECT 10.725 8.075 10.895 8.265 ;
        RECT 13.485 8.215 13.655 8.245 ;
        RECT 13.480 8.105 13.655 8.215 ;
        RECT 13.485 8.055 13.655 8.105 ;
        RECT 15.705 8.055 15.875 8.265 ;
        RECT 0.005 7.245 1.375 8.055 ;
        RECT 1.385 7.245 4.135 8.055 ;
        RECT 4.145 7.245 9.655 8.055 ;
        RECT 9.665 7.245 12.415 8.055 ;
        RECT 12.425 7.245 13.795 8.055 ;
        RECT 14.645 7.245 16.015 8.055 ;
        RECT 0.005 2.825 1.375 3.635 ;
        RECT 14.645 2.825 16.015 3.635 ;
        RECT 0.145 2.635 0.315 2.825 ;
        RECT 1.520 2.665 1.640 2.775 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 10.720 2.665 10.840 2.775 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 15.705 2.635 15.875 2.825 ;
      LAYER li1 ;
        RECT 1.925 2.975 2.445 4.460 ;
        RECT 3.305 2.975 3.825 4.460 ;
        RECT 4.685 2.975 5.205 4.460 ;
        RECT 6.065 2.975 6.585 4.460 ;
        RECT 7.445 2.975 7.965 4.460 ;
        RECT 8.825 2.975 9.345 4.460 ;
        RECT 11.125 2.975 11.645 4.460 ;
        RECT 12.505 2.975 13.025 4.460 ;
  END
END product_id_rom_8bit
END LIBRARY

