VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_routes
  CLASS COVER ;
  FOREIGN analog_routes ;
  ORIGIN 0.000 0.000 ;
  SIZE 3178.000 BY 4777.500 ;
  OBS
      LAYER met2 ;
        RECT 196.805 4778.265 198.375 4780.435 ;
        RECT 316.805 4778.265 318.375 4780.435 ;
        RECT 436.805 4778.265 438.375 4780.435 ;
        RECT 556.805 4778.265 558.375 4780.435 ;
        RECT 906.805 4778.265 908.375 4780.435 ;
        RECT 1026.805 4778.265 1028.375 4780.435 ;
        RECT 1146.805 4778.265 1148.375 4780.435 ;
        RECT 1266.805 4778.265 1268.375 4780.435 ;
        RECT 1481.805 4778.265 1483.375 4780.435 ;
        RECT 1596.805 4778.265 1598.375 4780.435 ;
        RECT 1636.310 4778.000 1638.120 4779.695 ;
        RECT 1639.400 4778.000 1642.655 4779.695 ;
        RECT 1961.805 4778.265 1963.375 4780.435 ;
        RECT 2081.805 4778.265 2083.375 4780.435 ;
        RECT 2201.805 4778.265 2203.375 4780.435 ;
        RECT 2321.805 4778.265 2323.375 4780.435 ;
        RECT 2671.805 4778.265 2673.375 4780.435 ;
        RECT 2791.805 4778.265 2793.375 4780.435 ;
        RECT 2911.805 4778.265 2913.375 4780.435 ;
        RECT 3031.805 4778.265 3033.375 4780.435 ;
        RECT 2677.665 50.220 2678.970 52.190 ;
        RECT 2679.830 50.215 2681.135 52.185 ;
        RECT 2724.750 50.135 2726.055 52.105 ;
        RECT 2841.245 49.620 2842.580 51.720 ;
        RECT 3058.895 49.615 3060.235 52.390 ;
      LAYER met3 ;
        RECT 196.655 4778.060 198.905 4780.435 ;
        RECT 316.655 4778.060 318.905 4780.435 ;
        RECT 436.655 4778.060 438.905 4780.435 ;
        RECT 556.655 4778.060 558.905 4780.435 ;
        RECT 906.655 4778.060 908.905 4780.435 ;
        RECT 1026.655 4778.060 1028.905 4780.435 ;
        RECT 1146.655 4778.060 1148.905 4780.435 ;
        RECT 1266.655 4778.060 1268.905 4780.435 ;
        RECT 1481.655 4778.060 1483.905 4780.435 ;
        RECT 1596.655 4778.060 1598.905 4780.435 ;
        RECT 1636.310 4778.000 1638.655 4779.695 ;
        RECT 1640.310 4778.000 1642.655 4779.695 ;
        RECT 1961.655 4778.060 1963.905 4780.435 ;
        RECT 2081.655 4778.060 2083.905 4780.435 ;
        RECT 2201.655 4778.060 2203.905 4780.435 ;
        RECT 2321.655 4778.060 2323.905 4780.435 ;
        RECT 2671.655 4778.060 2673.905 4780.435 ;
        RECT 2791.655 4778.060 2793.905 4780.435 ;
        RECT 2911.655 4778.060 2913.905 4780.435 ;
        RECT 3031.655 4778.060 3033.905 4780.435 ;
        RECT 3031.795 4777.430 3033.765 4778.060 ;
        RECT -2.370 4510.240 -0.110 4511.310 ;
        RECT 3178.425 4430.130 3180.685 4431.200 ;
        RECT -2.370 4405.240 -0.110 4406.310 ;
        RECT 3178.425 4325.140 3180.685 4326.210 ;
        RECT -2.370 4300.240 -0.110 4301.310 ;
        RECT 3178.425 4220.140 3180.685 4221.210 ;
        RECT -2.370 4195.240 -0.110 4196.310 ;
        RECT 3178.425 4115.140 3180.685 4116.210 ;
        RECT -2.290 3990.450 1.210 3991.090 ;
        RECT 3176.460 3909.915 3180.290 3910.560 ;
        RECT -2.290 3885.450 1.210 3886.090 ;
        RECT 3176.460 3804.915 3180.290 3805.560 ;
        RECT -2.290 3780.450 1.210 3781.090 ;
        RECT 3176.460 3699.915 3180.290 3700.560 ;
        RECT -2.290 3675.450 1.210 3676.090 ;
        RECT 3176.460 3594.915 3180.290 3595.560 ;
        RECT 3176.460 3144.405 3180.290 3144.450 ;
        RECT 3176.460 3143.805 3181.500 3144.405 ;
        RECT -2.290 3022.200 1.210 3022.240 ;
        RECT -3.500 3021.600 1.210 3022.200 ;
        RECT 3176.460 2979.405 3180.290 2979.450 ;
        RECT 3176.460 2978.805 3181.500 2979.405 ;
        RECT -2.290 2857.200 1.210 2857.240 ;
        RECT -3.500 2856.600 1.210 2857.200 ;
        RECT 3176.460 2814.405 3180.290 2814.450 ;
        RECT 3176.460 2813.805 3181.500 2814.405 ;
        RECT -2.290 2692.200 1.210 2692.240 ;
        RECT -3.500 2691.600 1.210 2692.200 ;
        RECT 3176.460 2649.405 3180.290 2649.450 ;
        RECT 3176.460 2648.805 3181.500 2649.405 ;
        RECT -2.290 2527.200 1.210 2527.240 ;
        RECT -3.500 2526.600 1.210 2527.200 ;
        RECT -0.645 2391.475 0.855 2391.620 ;
        RECT -2.185 2389.475 0.855 2391.475 ;
        RECT -0.645 2387.490 0.855 2389.475 ;
        RECT 3175.945 2377.805 3177.445 2378.020 ;
        RECT 3175.945 2375.805 3180.175 2377.805 ;
        RECT 3175.945 2373.890 3177.445 2375.805 ;
        RECT -2.290 2339.485 1.210 2340.125 ;
        RECT 3176.460 2330.480 3180.290 2330.525 ;
        RECT 3176.460 2329.880 3181.500 2330.480 ;
        RECT 3176.460 2161.405 3180.290 2161.450 ;
        RECT 3176.460 2160.805 3181.500 2161.405 ;
        RECT -2.290 2039.200 1.210 2039.240 ;
        RECT -2.295 2038.600 1.210 2039.200 ;
        RECT 3176.460 1996.405 3180.290 1996.450 ;
        RECT 3176.460 1995.805 3181.500 1996.405 ;
        RECT -2.290 1874.200 1.210 1874.240 ;
        RECT -3.500 1873.600 1.210 1874.200 ;
        RECT 3176.460 1830.120 3180.290 1830.165 ;
        RECT 3176.460 1829.520 3181.500 1830.120 ;
        RECT -2.290 1710.485 1.210 1710.525 ;
        RECT -3.500 1709.885 1.210 1710.485 ;
        RECT 3176.460 1665.120 3180.290 1665.165 ;
        RECT 3176.460 1664.520 3181.500 1665.120 ;
        RECT -2.290 1545.485 1.210 1545.525 ;
        RECT -3.500 1544.885 1.210 1545.485 ;
        RECT 2677.665 50.220 2678.970 52.190 ;
        RECT 2679.830 50.215 2681.135 52.185 ;
        RECT 2724.750 50.135 2726.055 52.105 ;
        RECT 2840.705 49.615 2842.580 52.685 ;
        RECT 3058.355 49.615 3060.230 52.685 ;
      LAYER met4 ;
        RECT 2998.185 4782.090 3001.385 4782.760 ;
        RECT 2998.095 4781.160 3001.385 4782.090 ;
        RECT 196.655 4778.060 198.905 4780.435 ;
        RECT 316.655 4778.060 318.905 4780.435 ;
        RECT 436.655 4778.060 438.905 4780.435 ;
        RECT 556.655 4778.060 558.905 4780.435 ;
        RECT 906.655 4778.060 908.905 4780.435 ;
        RECT 1026.655 4778.060 1028.905 4780.435 ;
        RECT 1146.655 4778.060 1148.905 4780.435 ;
        RECT 1266.655 4778.060 1268.905 4780.435 ;
        RECT 1481.655 4778.060 1483.905 4780.435 ;
        RECT 1596.655 4778.060 1598.905 4780.435 ;
        RECT 193.655 4629.595 194.655 4776.925 ;
        RECT 193.655 4625.595 195.255 4629.595 ;
        RECT 196.655 4624.850 197.655 4778.060 ;
        RECT 199.655 4629.595 200.655 4776.950 ;
        RECT 199.055 4625.595 200.655 4629.595 ;
        RECT 313.655 4629.595 314.655 4776.925 ;
        RECT 313.655 4625.595 315.255 4629.595 ;
        RECT 316.655 4624.850 317.655 4778.060 ;
        RECT 319.655 4629.595 320.655 4776.950 ;
        RECT 319.055 4625.595 320.655 4629.595 ;
        RECT 433.655 4629.595 434.655 4776.925 ;
        RECT 433.655 4625.595 435.255 4629.595 ;
        RECT 436.655 4624.850 437.655 4778.060 ;
        RECT 439.655 4629.595 440.655 4776.950 ;
        RECT 439.055 4625.595 440.655 4629.595 ;
        RECT 553.655 4629.595 554.655 4776.925 ;
        RECT 553.655 4625.595 555.255 4629.595 ;
        RECT 556.655 4624.850 557.655 4778.060 ;
        RECT 559.655 4629.595 560.655 4776.950 ;
        RECT 559.055 4625.595 560.655 4629.595 ;
        RECT 903.655 4629.595 904.655 4776.925 ;
        RECT 903.655 4625.595 905.255 4629.595 ;
        RECT 906.655 4624.850 907.655 4778.060 ;
        RECT 909.655 4629.595 910.655 4776.950 ;
        RECT 909.055 4625.595 910.655 4629.595 ;
        RECT 1023.655 4629.595 1024.655 4776.925 ;
        RECT 1023.655 4625.595 1025.255 4629.595 ;
        RECT 1026.655 4624.850 1027.655 4778.060 ;
        RECT 1029.655 4629.595 1030.655 4776.950 ;
        RECT 1029.055 4625.595 1030.655 4629.595 ;
        RECT 1143.655 4629.595 1144.655 4776.925 ;
        RECT 1143.655 4625.595 1145.255 4629.595 ;
        RECT 1146.655 4624.850 1147.655 4778.060 ;
        RECT 1149.655 4629.595 1150.655 4776.950 ;
        RECT 1149.055 4625.595 1150.655 4629.595 ;
        RECT 1263.655 4629.595 1264.655 4776.925 ;
        RECT 1263.655 4625.595 1265.255 4629.595 ;
        RECT 1266.655 4624.850 1267.655 4778.060 ;
        RECT 1269.655 4629.595 1270.655 4776.950 ;
        RECT 1269.055 4625.595 1270.655 4629.595 ;
        RECT 1478.655 4629.595 1479.655 4776.925 ;
        RECT 1478.655 4625.595 1480.255 4629.595 ;
        RECT 1481.655 4624.850 1482.655 4778.060 ;
        RECT 1484.655 4629.595 1485.655 4776.950 ;
        RECT 1484.055 4625.595 1485.655 4629.595 ;
        RECT 1593.655 4629.595 1594.655 4776.925 ;
        RECT 1593.655 4625.595 1595.255 4629.595 ;
        RECT 1596.655 4624.850 1597.655 4778.060 ;
        RECT 1636.310 4778.000 1638.655 4779.695 ;
        RECT 1640.310 4778.000 1642.655 4779.695 ;
        RECT 1599.655 4629.595 1600.655 4776.950 ;
        RECT 1599.055 4625.595 1600.655 4629.595 ;
        RECT 1635.655 4624.850 1636.655 4777.080 ;
        RECT 1637.655 4624.850 1638.655 4778.000 ;
        RECT 1639.655 4624.850 1640.655 4777.080 ;
        RECT 1641.655 4624.850 1642.655 4778.000 ;
        RECT 1961.655 4778.060 1963.905 4780.435 ;
        RECT 2081.655 4778.060 2083.905 4780.435 ;
        RECT 2201.655 4778.060 2203.905 4780.435 ;
        RECT 2321.655 4778.060 2323.905 4780.435 ;
        RECT 2671.655 4778.060 2673.905 4780.435 ;
        RECT 2791.655 4778.060 2793.905 4780.435 ;
        RECT 2911.655 4778.060 2913.905 4780.435 ;
        RECT 1643.655 4624.850 1644.655 4777.080 ;
        RECT 1958.655 4629.595 1959.655 4776.925 ;
        RECT 1958.655 4625.595 1960.255 4629.595 ;
        RECT 1961.655 4624.850 1962.655 4778.060 ;
        RECT 1964.655 4629.595 1965.655 4776.950 ;
        RECT 1964.055 4625.595 1965.655 4629.595 ;
        RECT 2078.655 4629.595 2079.655 4776.925 ;
        RECT 2078.655 4625.595 2080.255 4629.595 ;
        RECT 2081.655 4624.850 2082.655 4778.060 ;
        RECT 2084.655 4629.595 2085.655 4776.950 ;
        RECT 2084.055 4625.595 2085.655 4629.595 ;
        RECT 2198.655 4629.595 2199.655 4776.925 ;
        RECT 2198.655 4625.595 2200.255 4629.595 ;
        RECT 2201.655 4624.850 2202.655 4778.060 ;
        RECT 2204.655 4629.595 2205.655 4776.950 ;
        RECT 2204.055 4625.595 2205.655 4629.595 ;
        RECT 2318.655 4629.595 2319.655 4776.925 ;
        RECT 2318.655 4625.595 2320.255 4629.595 ;
        RECT 2321.655 4624.850 2322.655 4778.060 ;
        RECT 2324.655 4629.595 2325.655 4776.950 ;
        RECT 2324.055 4625.595 2325.655 4629.595 ;
        RECT 2668.655 4629.595 2669.655 4776.925 ;
        RECT 2668.655 4625.595 2670.255 4629.595 ;
        RECT 2671.655 4624.850 2672.655 4778.060 ;
        RECT 2674.655 4629.595 2675.655 4776.950 ;
        RECT 2674.055 4625.595 2675.655 4629.595 ;
        RECT 2788.655 4629.595 2789.655 4776.925 ;
        RECT 2788.655 4625.595 2790.255 4629.595 ;
        RECT 2791.655 4624.850 2792.655 4778.060 ;
        RECT 2794.655 4629.595 2795.655 4776.950 ;
        RECT 2794.055 4625.595 2795.655 4629.595 ;
        RECT 2908.655 4629.595 2909.655 4776.925 ;
        RECT 2908.655 4625.595 2910.255 4629.595 ;
        RECT 2911.655 4624.850 2912.655 4778.060 ;
        RECT 2914.655 4629.595 2915.655 4776.950 ;
        RECT 2914.055 4625.595 2915.655 4629.595 ;
        RECT 2998.095 4629.595 2999.095 4781.160 ;
        RECT 3031.655 4779.390 3033.905 4779.635 ;
        RECT 3001.215 4778.680 3004.415 4779.210 ;
        RECT 3001.095 4777.610 3004.415 4778.680 ;
        RECT 3030.565 4777.790 3033.905 4779.390 ;
        RECT 2998.095 4625.595 2999.695 4629.595 ;
        RECT 3001.095 4624.850 3002.095 4777.610 ;
        RECT 3031.655 4777.260 3033.905 4777.790 ;
        RECT 3004.195 4775.100 3007.395 4775.720 ;
        RECT 3004.095 4774.120 3007.395 4775.100 ;
        RECT 3004.095 4629.595 3005.095 4774.120 ;
        RECT 3003.495 4625.595 3005.095 4629.595 ;
        RECT -2.535 4509.950 3.230 4511.550 ;
        RECT 146.490 4504.950 151.490 4516.560 ;
        RECT 3026.825 4424.840 3031.825 4436.450 ;
        RECT 3175.085 4429.840 3180.850 4431.440 ;
        RECT -2.535 4404.950 3.230 4406.550 ;
        RECT 146.490 4399.950 151.490 4411.560 ;
        RECT 3026.825 4319.850 3031.825 4331.460 ;
        RECT 3175.085 4324.850 3180.850 4326.450 ;
        RECT -2.535 4299.950 3.230 4301.550 ;
        RECT 146.490 4294.950 151.490 4306.560 ;
        RECT 3026.825 4214.850 3031.825 4226.460 ;
        RECT 3175.085 4219.850 3180.850 4221.450 ;
        RECT -2.535 4194.950 3.230 4196.550 ;
        RECT 146.490 4189.950 151.490 4201.560 ;
        RECT 3026.825 4109.850 3031.825 4121.460 ;
        RECT 3175.085 4114.850 3180.850 4116.450 ;
        RECT 153.135 3996.630 153.775 4048.850 ;
        RECT 150.570 3995.030 153.775 3996.630 ;
        RECT 153.135 3995.025 153.775 3995.030 ;
        RECT 154.435 3991.630 155.075 4048.850 ;
        RECT -1.240 3991.090 1.240 3991.630 ;
        RECT -2.290 3990.450 1.240 3991.090 ;
        RECT -1.240 3990.030 1.240 3990.450 ;
        RECT 151.875 3990.030 155.075 3991.630 ;
        RECT 155.695 3986.630 156.335 4048.850 ;
        RECT 153.135 3985.030 156.335 3986.630 ;
        RECT 155.695 3891.630 156.335 3985.030 ;
        RECT 153.130 3890.030 156.335 3891.630 ;
        RECT 155.695 3890.020 156.335 3890.030 ;
        RECT 156.995 3886.630 157.635 4048.850 ;
        RECT -1.240 3886.090 1.240 3886.630 ;
        RECT -2.290 3885.450 1.240 3886.090 ;
        RECT -1.240 3885.030 1.240 3885.450 ;
        RECT 154.440 3885.030 157.640 3886.630 ;
        RECT 158.255 3881.630 158.895 4048.850 ;
        RECT 155.695 3880.030 158.895 3881.630 ;
        RECT 158.255 3786.635 158.895 3880.030 ;
        RECT 155.695 3785.035 158.895 3786.635 ;
        RECT 158.255 3785.025 158.895 3785.035 ;
        RECT 159.555 3781.630 160.195 4048.850 ;
        RECT -1.240 3781.090 1.240 3781.630 ;
        RECT -2.290 3780.450 1.240 3781.090 ;
        RECT -1.240 3780.030 1.240 3780.450 ;
        RECT 156.995 3780.030 160.195 3781.630 ;
        RECT 160.815 3776.625 161.455 4048.850 ;
        RECT 158.250 3775.025 161.455 3776.625 ;
        RECT 160.815 3681.630 161.455 3775.025 ;
        RECT 158.255 3680.030 161.455 3681.630 ;
        RECT 160.815 3679.980 161.455 3680.030 ;
        RECT 162.115 3676.630 162.755 4048.850 ;
        RECT -1.240 3676.090 1.240 3676.630 ;
        RECT -2.290 3675.450 1.240 3676.090 ;
        RECT -1.240 3675.030 1.240 3675.450 ;
        RECT 159.560 3675.030 162.760 3676.630 ;
        RECT 163.375 3671.640 164.015 4048.850 ;
        RECT 160.820 3670.040 164.020 3671.640 ;
        RECT 163.375 3027.770 164.015 3670.040 ;
        RECT 160.815 3026.170 164.015 3027.770 ;
        RECT 164.675 3022.790 165.315 4048.850 ;
        RECT -1.240 3022.240 1.240 3022.785 ;
        RECT -2.290 3021.600 1.240 3022.240 ;
        RECT -1.240 3021.180 1.240 3021.600 ;
        RECT 162.115 3021.190 165.315 3022.790 ;
        RECT 165.935 3017.770 166.575 4048.850 ;
        RECT 163.380 3016.170 166.580 3017.770 ;
        RECT 165.935 2862.765 166.575 3016.170 ;
        RECT 163.380 2861.165 166.580 2862.765 ;
        RECT 165.935 2861.145 166.575 2861.165 ;
        RECT -1.240 2857.240 1.240 2857.780 ;
        RECT 167.235 2857.760 167.875 4048.850 ;
        RECT -2.290 2856.600 1.240 2857.240 ;
        RECT -1.240 2856.180 1.240 2856.600 ;
        RECT 164.675 2856.160 167.875 2857.760 ;
        RECT 168.495 2852.770 169.135 4048.850 ;
        RECT 165.935 2851.170 169.135 2852.770 ;
        RECT 168.495 2697.890 169.135 2851.170 ;
        RECT 165.940 2696.290 169.140 2697.890 ;
        RECT 168.495 2696.270 169.135 2696.290 ;
        RECT 169.795 2692.900 170.435 4048.850 ;
        RECT -1.240 2692.240 1.240 2692.780 ;
        RECT -2.290 2691.600 1.240 2692.240 ;
        RECT -1.240 2691.180 1.240 2691.600 ;
        RECT 167.235 2691.300 170.435 2692.900 ;
        RECT 171.055 2687.905 171.695 4048.850 ;
        RECT 168.500 2686.305 171.700 2687.905 ;
        RECT 171.055 2532.765 171.695 2686.305 ;
        RECT 168.495 2531.165 171.695 2532.765 ;
        RECT -1.240 2527.240 1.240 2527.780 ;
        RECT 172.355 2527.775 172.995 4048.850 ;
        RECT -2.290 2526.600 1.240 2527.240 ;
        RECT -1.240 2526.180 1.240 2526.600 ;
        RECT 169.795 2526.175 172.995 2527.775 ;
        RECT 173.615 2522.770 174.255 4048.850 ;
        RECT 171.065 2521.170 174.265 2522.770 ;
        RECT -0.645 2387.490 0.855 2391.620 ;
        RECT -0.275 2340.665 0.485 2387.490 ;
        RECT 173.615 2345.670 174.255 2521.170 ;
        RECT 171.055 2344.070 174.255 2345.670 ;
        RECT 173.615 2344.060 174.255 2344.070 ;
        RECT 174.915 2340.665 175.555 4048.850 ;
        RECT -1.240 2340.125 1.240 2340.665 ;
        RECT -2.290 2339.485 1.240 2340.125 ;
        RECT -1.240 2339.065 1.240 2339.485 ;
        RECT 172.355 2339.065 175.555 2340.665 ;
        RECT 176.175 2335.670 176.815 4048.850 ;
        RECT 173.610 2334.070 176.815 2335.670 ;
        RECT 176.175 2044.765 176.815 2334.070 ;
        RECT 173.615 2043.165 176.815 2044.765 ;
        RECT -1.240 2039.240 1.240 2039.780 ;
        RECT 177.475 2039.775 178.115 4048.850 ;
        RECT -2.290 2038.600 1.240 2039.240 ;
        RECT -1.240 2038.180 1.240 2038.600 ;
        RECT 174.925 2038.175 178.125 2039.775 ;
        RECT 178.735 2034.775 179.375 4048.850 ;
        RECT 176.175 2033.175 179.375 2034.775 ;
        RECT 178.735 1879.760 179.375 2033.175 ;
        RECT 176.165 1878.170 179.375 1879.760 ;
        RECT 176.165 1878.160 179.365 1878.170 ;
        RECT -1.240 1874.240 1.240 1874.780 ;
        RECT 180.035 1874.760 180.675 4048.850 ;
        RECT -2.290 1873.600 1.240 1874.240 ;
        RECT -1.240 1873.180 1.240 1873.600 ;
        RECT 177.475 1873.160 180.675 1874.760 ;
        RECT 181.295 1869.760 181.935 4048.850 ;
        RECT 178.735 1868.160 181.935 1869.760 ;
        RECT 181.295 1716.070 181.935 1868.160 ;
        RECT 178.735 1714.470 181.935 1716.070 ;
        RECT -1.240 1710.525 1.240 1711.065 ;
        RECT 182.595 1711.040 183.235 4048.850 ;
        RECT -2.290 1709.885 1.240 1710.525 ;
        RECT -1.240 1709.465 1.240 1709.885 ;
        RECT 180.035 1709.440 183.235 1711.040 ;
        RECT 183.855 1706.070 184.495 4048.850 ;
        RECT 181.300 1704.470 184.500 1706.070 ;
        RECT 183.855 1551.040 184.495 1704.470 ;
        RECT 181.175 1549.440 184.495 1551.040 ;
        RECT 183.855 1549.400 184.495 1549.440 ;
        RECT -1.240 1545.525 1.240 1546.065 ;
        RECT 185.155 1546.060 185.795 4048.850 ;
        RECT -2.290 1544.885 1.240 1545.525 ;
        RECT -1.240 1544.465 1.240 1544.885 ;
        RECT 182.595 1544.460 185.795 1546.060 ;
        RECT 186.455 1541.185 187.095 4048.850 ;
        RECT 1882.595 3851.060 1883.235 4048.850 ;
        RECT 1883.875 3848.850 1884.515 4048.850 ;
        RECT 1885.155 3851.060 1885.795 4048.850 ;
        RECT 1886.435 3848.850 1887.075 4048.850 ;
        RECT 1887.715 3851.060 1888.355 4048.850 ;
        RECT 1888.995 3848.850 1889.635 4048.850 ;
        RECT 1890.275 3851.060 1890.915 4048.850 ;
        RECT 1891.555 3848.850 1892.195 4048.850 ;
        RECT 1892.835 3851.060 1893.475 4048.850 ;
        RECT 1894.115 3848.850 1894.755 4048.850 ;
        RECT 1895.395 3851.060 1896.035 4048.850 ;
        RECT 1896.675 3848.850 1897.315 4048.850 ;
        RECT 1897.955 3851.060 1898.595 4048.850 ;
        RECT 1899.235 3848.850 1899.875 4048.850 ;
        RECT 1900.515 3851.060 1901.155 4048.850 ;
        RECT 1901.795 3848.850 1902.435 4048.850 ;
        RECT 1903.075 3851.060 1903.715 4048.850 ;
        RECT 1904.355 3848.850 1904.995 4048.850 ;
        RECT 1905.635 3851.060 1906.275 4048.850 ;
        RECT 1906.915 3848.850 1907.555 4048.850 ;
        RECT 1908.195 3851.060 1908.835 4048.850 ;
        RECT 1909.475 3848.850 1910.115 4048.850 ;
        RECT 1910.755 3851.060 1911.395 4048.850 ;
        RECT 1912.035 3848.850 1912.675 4048.850 ;
        RECT 1913.315 3851.060 1913.955 4048.850 ;
        RECT 1914.595 3848.850 1915.235 4048.850 ;
        RECT 1915.875 3851.060 1916.515 4048.850 ;
        RECT 1917.155 3848.850 1917.795 4048.850 ;
        RECT 1918.435 3851.060 1919.075 4048.850 ;
        RECT 1919.715 3848.850 1920.355 4048.850 ;
        RECT 1920.995 3851.060 1921.635 4048.850 ;
        RECT 1922.275 3848.850 1922.915 4048.850 ;
        RECT 1923.555 3851.060 1924.195 4048.850 ;
        RECT 1924.835 3848.850 1925.475 4048.850 ;
        RECT 1926.115 3851.060 1926.755 4048.850 ;
        RECT 1927.395 3848.850 1928.035 4048.850 ;
        RECT 1928.675 3851.060 1929.315 4048.850 ;
        RECT 1929.955 3848.850 1930.595 4048.850 ;
        RECT 1931.235 3851.060 1931.875 4048.850 ;
        RECT 1932.515 3848.850 1933.155 4048.850 ;
        RECT 1933.795 3851.060 1934.435 4048.850 ;
        RECT 1935.075 3848.850 1935.715 4048.850 ;
        RECT 1936.355 3851.060 1936.995 4048.850 ;
        RECT 1937.635 3848.850 1938.275 4048.850 ;
        RECT 1938.915 3851.060 1939.555 4048.850 ;
        RECT 1940.195 3848.850 1940.835 4048.850 ;
        RECT 1941.475 3851.060 1942.115 4048.850 ;
        RECT 1942.755 3848.850 1943.395 4048.850 ;
        RECT 1944.035 3851.060 1944.675 4048.850 ;
        RECT 1945.315 3848.850 1945.955 4048.850 ;
        RECT 1946.595 3851.060 1947.235 4048.850 ;
        RECT 1947.875 3848.850 1948.515 4048.850 ;
        RECT 1949.155 3851.060 1949.795 4048.850 ;
        RECT 1950.435 3848.850 1951.075 4048.850 ;
        RECT 1951.715 3851.060 1952.355 4048.850 ;
        RECT 1952.995 3848.850 1953.635 4048.850 ;
        RECT 1954.275 3851.060 1954.915 4048.850 ;
        RECT 1955.555 3848.850 1956.195 4048.850 ;
        RECT 1956.835 3851.060 1957.475 4048.850 ;
        RECT 1958.115 3848.850 1958.755 4048.850 ;
        RECT 1959.395 3851.060 1960.035 4048.850 ;
        RECT 1960.675 3848.850 1961.315 4048.850 ;
        RECT 1961.955 3851.070 1962.595 4048.850 ;
        RECT 1963.235 3848.850 1963.875 4048.850 ;
        RECT 1964.515 3851.060 1965.155 4048.850 ;
        RECT 1965.795 3848.850 1966.435 4048.850 ;
        RECT 1967.075 3851.070 1967.715 4048.850 ;
        RECT 2963.375 1635.090 2964.015 4048.855 ;
        RECT 2964.675 1636.390 2965.315 4048.855 ;
        RECT 2965.935 1637.650 2966.575 4048.855 ;
        RECT 2967.235 1638.950 2967.875 4048.855 ;
        RECT 2968.495 1640.210 2969.135 4048.855 ;
        RECT 2969.795 1641.510 2970.435 4048.855 ;
        RECT 2971.055 1642.770 2971.695 4048.855 ;
        RECT 2972.355 1644.070 2972.995 4048.855 ;
        RECT 2973.615 1645.330 2974.255 4048.855 ;
        RECT 2974.915 1646.630 2975.555 4048.855 ;
        RECT 2976.175 1647.890 2976.815 4048.855 ;
        RECT 2977.475 1649.190 2978.115 4048.855 ;
        RECT 2978.735 1650.450 2979.375 4048.855 ;
        RECT 2980.035 1651.750 2980.675 4048.855 ;
        RECT 2981.295 1660.680 2981.935 4048.855 ;
        RECT 2982.595 1665.670 2983.235 4048.855 ;
        RECT 2983.895 1825.540 2984.535 4048.855 ;
        RECT 2985.155 1830.525 2985.795 4048.855 ;
        RECT 2986.455 1991.905 2987.095 4048.855 ;
        RECT 2987.715 1996.965 2988.355 4048.855 ;
        RECT 2989.015 2157.000 2989.655 4048.855 ;
        RECT 2990.275 2161.970 2990.915 4048.855 ;
        RECT 2991.575 2325.985 2992.215 4048.855 ;
        RECT 2992.835 2331.030 2993.475 4048.855 ;
        RECT 2994.135 2644.960 2994.775 4048.855 ;
        RECT 2995.395 2649.970 2996.035 4048.855 ;
        RECT 2996.695 2809.910 2997.335 4048.855 ;
        RECT 2997.955 2814.970 2998.595 4048.855 ;
        RECT 2999.255 2974.975 2999.895 4048.855 ;
        RECT 3000.515 2979.970 3001.155 4048.855 ;
        RECT 3001.815 3140.065 3002.455 4048.855 ;
        RECT 3003.075 3144.975 3003.715 4048.855 ;
        RECT 3004.375 3591.020 3005.015 4048.855 ;
        RECT 3005.635 3596.065 3006.275 4048.855 ;
        RECT 3006.935 3696.040 3007.575 4048.855 ;
        RECT 3008.195 3701.095 3008.835 4048.855 ;
        RECT 3009.495 3801.025 3010.135 4048.855 ;
        RECT 3010.755 3806.145 3011.395 4048.855 ;
        RECT 3012.055 3906.075 3012.695 4048.855 ;
        RECT 3013.315 3911.065 3013.955 4048.855 ;
        RECT 3014.615 3916.070 3015.255 4048.855 ;
        RECT 3014.615 3914.810 3017.890 3916.070 ;
        RECT 3014.690 3914.470 3017.890 3914.810 ;
        RECT 3013.310 3909.465 3016.510 3911.065 ;
        RECT 3175.160 3910.560 3178.605 3911.065 ;
        RECT 3175.160 3909.915 3180.290 3910.560 ;
        RECT 3175.160 3909.465 3178.605 3909.915 ;
        RECT 3012.055 3904.475 3015.305 3906.075 ;
        RECT 3012.055 3811.030 3012.695 3904.475 ;
        RECT 3012.020 3809.430 3015.220 3811.030 ;
        RECT 3010.750 3804.545 3013.950 3806.145 ;
        RECT 3175.160 3805.560 3178.605 3806.065 ;
        RECT 3175.160 3804.915 3180.290 3805.560 ;
        RECT 3175.160 3804.465 3178.605 3804.915 ;
        RECT 3009.495 3799.425 3012.730 3801.025 ;
        RECT 3009.495 3706.015 3010.135 3799.425 ;
        RECT 3009.495 3704.415 3012.705 3706.015 ;
        RECT 3009.495 3704.170 3010.135 3704.415 ;
        RECT 3008.190 3699.495 3011.390 3701.095 ;
        RECT 3175.160 3700.560 3178.605 3701.065 ;
        RECT 3175.160 3699.915 3180.290 3700.560 ;
        RECT 3175.160 3699.465 3178.605 3699.915 ;
        RECT 3006.935 3694.440 3010.245 3696.040 ;
        RECT 3006.935 3601.030 3007.575 3694.440 ;
        RECT 3006.935 3599.430 3010.165 3601.030 ;
        RECT 3006.935 3599.280 3007.575 3599.430 ;
        RECT 3005.455 3594.465 3008.655 3596.065 ;
        RECT 3175.160 3595.560 3178.605 3596.065 ;
        RECT 3175.160 3594.915 3180.290 3595.560 ;
        RECT 3175.160 3594.465 3178.605 3594.915 ;
        RECT 3004.375 3589.420 3007.615 3591.020 ;
        RECT 3004.375 3150.100 3005.015 3589.420 ;
        RECT 3004.375 3148.500 3007.585 3150.100 ;
        RECT 3004.375 3148.415 3005.015 3148.500 ;
        RECT 3003.070 3143.375 3006.270 3144.975 ;
        RECT 3175.160 3144.450 3178.605 3144.955 ;
        RECT 3175.160 3143.805 3180.290 3144.450 ;
        RECT 3175.160 3143.355 3178.605 3143.805 ;
        RECT 3001.815 3138.465 3005.025 3140.065 ;
        RECT 3001.815 2984.950 3002.455 3138.465 ;
        RECT 3001.815 2983.350 3005.135 2984.950 ;
        RECT 3001.815 2983.100 3002.455 2983.350 ;
        RECT 3000.335 2978.370 3003.535 2979.970 ;
        RECT 3175.160 2979.450 3178.605 2979.955 ;
        RECT 3175.160 2978.805 3180.290 2979.450 ;
        RECT 3175.160 2978.355 3178.605 2978.805 ;
        RECT 2999.250 2973.375 3002.450 2974.975 ;
        RECT 2999.255 2819.885 2999.895 2973.375 ;
        RECT 2999.220 2818.285 3002.420 2819.885 ;
        RECT 2997.775 2813.370 3000.975 2814.970 ;
        RECT 3175.160 2814.450 3178.605 2814.955 ;
        RECT 3175.160 2813.805 3180.290 2814.450 ;
        RECT 3175.160 2813.355 3178.605 2813.805 ;
        RECT 2996.685 2808.310 2999.885 2809.910 ;
        RECT 2996.695 2654.965 2997.335 2808.310 ;
        RECT 2996.695 2653.365 2999.915 2654.965 ;
        RECT 2996.695 2652.805 2997.335 2653.365 ;
        RECT 2995.215 2648.370 2998.415 2649.970 ;
        RECT 3175.160 2649.450 3178.605 2649.955 ;
        RECT 3175.160 2648.805 3180.290 2649.450 ;
        RECT 3175.160 2648.355 3178.605 2648.805 ;
        RECT 2994.135 2643.360 2997.345 2644.960 ;
        RECT 2994.135 2336.020 2994.775 2643.360 ;
        RECT 3176.345 2378.020 3177.105 2378.050 ;
        RECT 3175.945 2373.890 3177.445 2378.020 ;
        RECT 2994.135 2334.420 2997.345 2336.020 ;
        RECT 2994.135 2333.805 2994.775 2334.420 ;
        RECT 3176.345 2331.030 3177.105 2373.890 ;
        RECT 2992.655 2329.430 2995.855 2331.030 ;
        RECT 3175.160 2330.525 3178.605 2331.030 ;
        RECT 3175.160 2329.880 3180.290 2330.525 ;
        RECT 3175.160 2329.430 3178.605 2329.880 ;
        RECT 2991.550 2324.385 2994.750 2325.985 ;
        RECT 2991.575 2166.885 2992.215 2324.385 ;
        RECT 2991.550 2165.285 2994.750 2166.885 ;
        RECT 2991.575 2164.930 2992.215 2165.285 ;
        RECT 2990.095 2160.370 2993.295 2161.970 ;
        RECT 3175.160 2161.450 3178.605 2161.955 ;
        RECT 3175.160 2160.805 3180.290 2161.450 ;
        RECT 3175.160 2160.355 3178.605 2160.805 ;
        RECT 2989.015 2155.400 2992.270 2157.000 ;
        RECT 2989.015 2001.910 2989.655 2155.400 ;
        RECT 2989.010 2000.310 2992.210 2001.910 ;
        RECT 2989.015 2000.120 2989.655 2000.310 ;
        RECT 2987.535 1995.365 2990.735 1996.965 ;
        RECT 3175.160 1996.450 3178.605 1996.955 ;
        RECT 3175.160 1995.805 3180.290 1996.450 ;
        RECT 3175.160 1995.355 3178.605 1995.805 ;
        RECT 2986.455 1990.305 2989.760 1991.905 ;
        RECT 2986.455 1835.600 2987.095 1990.305 ;
        RECT 2986.385 1834.000 2989.585 1835.600 ;
        RECT 2985.025 1828.925 2988.225 1830.525 ;
        RECT 3175.160 1830.165 3178.605 1830.670 ;
        RECT 3175.160 1829.520 3180.290 1830.165 ;
        RECT 3175.160 1829.070 3178.605 1829.520 ;
        RECT 2983.895 1823.940 2987.135 1825.540 ;
        RECT 2983.895 1670.685 2984.535 1823.940 ;
        RECT 2983.880 1669.085 2987.080 1670.685 ;
        RECT 2982.465 1664.070 2985.665 1665.670 ;
        RECT 3175.160 1665.165 3178.605 1665.670 ;
        RECT 3175.160 1664.520 3180.290 1665.165 ;
        RECT 3175.160 1664.070 3178.605 1664.520 ;
        RECT 2981.280 1659.080 2984.480 1660.680 ;
        RECT 2981.295 1653.010 2981.935 1659.080 ;
        RECT 2981.295 1652.370 3031.935 1653.010 ;
        RECT 2980.035 1651.110 3030.675 1651.750 ;
        RECT 2978.735 1649.810 3029.375 1650.450 ;
        RECT 2977.475 1648.550 3028.115 1649.190 ;
        RECT 2976.175 1647.250 3026.815 1647.890 ;
        RECT 2974.915 1645.990 3025.555 1646.630 ;
        RECT 2973.615 1644.690 3024.255 1645.330 ;
        RECT 2972.355 1643.430 3022.995 1644.070 ;
        RECT 2971.055 1642.130 3021.695 1642.770 ;
        RECT 2969.795 1640.870 3020.435 1641.510 ;
        RECT 2968.495 1639.570 3019.135 1640.210 ;
        RECT 2967.235 1638.310 3017.875 1638.950 ;
        RECT 2965.935 1637.010 3016.575 1637.650 ;
        RECT 2964.675 1635.750 3015.315 1636.390 ;
        RECT 3013.375 1635.090 3014.015 1635.095 ;
        RECT 2963.375 1634.465 3014.015 1635.090 ;
        RECT 2992.070 1634.450 3014.015 1634.465 ;
        RECT 183.775 1539.585 187.095 1541.185 ;
        RECT 186.455 1539.465 187.095 1539.585 ;
        RECT 3013.375 109.320 3014.015 1634.450 ;
        RECT 2641.475 109.175 2644.675 109.290 ;
        RECT 2641.440 107.690 2644.675 109.175 ;
        RECT 3010.820 107.720 3014.020 109.320 ;
        RECT 2641.440 12.070 2643.040 107.690 ;
        RECT 2644.710 104.190 2646.610 104.370 ;
        RECT 3014.675 104.275 3015.315 1635.750 ;
        RECT 2644.710 102.590 2648.030 104.190 ;
        RECT 3012.070 103.585 3015.315 104.275 ;
        RECT 3012.070 102.675 3015.270 103.585 ;
        RECT 2644.710 102.470 2646.610 102.590 ;
        RECT 2639.880 10.470 2643.080 12.070 ;
        RECT 2644.940 8.715 2646.540 102.470 ;
        RECT 2648.535 98.820 2651.735 99.305 ;
        RECT 3015.935 99.295 3016.575 1637.010 ;
        RECT 2648.440 97.705 2651.735 98.820 ;
        RECT 3013.300 98.300 3016.575 99.295 ;
        RECT 2644.795 8.565 2646.695 8.715 ;
        RECT 2643.305 6.965 2646.695 8.565 ;
        RECT 2644.795 6.815 2646.695 6.965 ;
        RECT 2648.440 5.120 2650.040 97.705 ;
        RECT 3013.300 97.695 3016.500 98.300 ;
        RECT 2651.790 94.230 2653.690 94.410 ;
        RECT 3017.235 94.340 3017.875 1638.310 ;
        RECT 2651.790 92.630 2655.110 94.230 ;
        RECT 3014.530 93.485 3017.875 94.340 ;
        RECT 3014.530 92.740 3017.730 93.485 ;
        RECT 2651.790 92.510 2653.690 92.630 ;
        RECT 2646.815 3.665 2650.040 5.120 ;
        RECT 2646.815 3.520 2650.015 3.665 ;
        RECT 2651.940 1.745 2653.540 92.510 ;
        RECT 2655.440 89.250 2657.040 89.630 ;
        RECT 3018.495 89.275 3019.135 1639.570 ;
        RECT 2655.440 87.650 2658.765 89.250 ;
        RECT 3015.865 88.280 3019.135 89.275 ;
        RECT 3015.865 87.675 3019.065 88.280 ;
        RECT 2651.695 1.675 2653.595 1.745 ;
        RECT 2650.240 0.075 2653.595 1.675 ;
        RECT 2651.695 -0.155 2653.595 0.075 ;
        RECT 2655.440 -1.770 2657.040 87.650 ;
        RECT 2677.440 84.400 2679.220 84.405 ;
        RECT 2677.385 84.220 2679.285 84.400 ;
        RECT 3019.795 84.325 3020.435 1640.870 ;
        RECT 2677.385 82.620 2680.705 84.220 ;
        RECT 3017.115 84.110 3020.435 84.325 ;
        RECT 3017.115 82.725 3020.315 84.110 ;
        RECT 2677.385 82.500 2679.285 82.620 ;
        RECT 2677.605 50.165 2679.030 82.500 ;
        RECT 3021.055 79.360 3021.695 1642.130 ;
        RECT 3018.425 77.760 3021.695 79.360 ;
        RECT 3021.055 77.555 3021.695 77.760 ;
        RECT 2679.540 74.250 2681.440 74.430 ;
        RECT 3022.355 74.375 3022.995 1643.430 ;
        RECT 2679.540 72.650 2682.860 74.250 ;
        RECT 3019.715 72.775 3022.995 74.375 ;
        RECT 2679.540 72.530 2681.440 72.650 ;
        RECT 3022.355 72.635 3022.995 72.775 ;
        RECT 2679.735 50.125 2681.180 72.530 ;
        RECT 3023.615 69.300 3024.255 1644.690 ;
        RECT 3020.920 68.400 3024.255 69.300 ;
        RECT 3020.920 67.700 3024.120 68.400 ;
        RECT 2724.440 64.215 2726.340 64.395 ;
        RECT 3024.915 64.335 3025.555 1645.990 ;
        RECT 2724.440 62.615 2727.760 64.215 ;
        RECT 3022.210 64.205 3025.555 64.335 ;
        RECT 3022.210 62.735 3025.410 64.205 ;
        RECT 2724.440 62.495 2726.340 62.615 ;
        RECT 2724.655 50.050 2726.155 62.495 ;
        RECT 3026.175 59.305 3026.815 1647.250 ;
        RECT 3023.480 57.705 3026.815 59.305 ;
        RECT 3026.175 57.630 3026.815 57.705 ;
        RECT 2840.710 54.355 2842.580 54.525 ;
        RECT 3027.475 54.405 3028.115 1648.550 ;
        RECT 2840.690 54.255 2842.580 54.355 ;
        RECT 3024.860 54.300 3028.115 54.405 ;
        RECT 2840.690 52.670 2843.995 54.255 ;
        RECT 3024.860 52.805 3028.060 54.300 ;
        RECT 2840.710 52.655 2843.995 52.670 ;
        RECT 2840.710 49.620 2842.580 52.655 ;
        RECT 3028.735 49.405 3029.375 1649.810 ;
        RECT 3030.035 54.405 3030.675 1651.110 ;
        RECT 3031.295 59.205 3031.935 1652.370 ;
        RECT 3031.295 57.605 3034.685 59.205 ;
        RECT 3031.295 57.355 3031.935 57.605 ;
        RECT 3030.035 54.305 3033.305 54.405 ;
        RECT 3030.105 52.805 3033.305 54.305 ;
        RECT 3058.360 54.255 3060.230 54.295 ;
        RECT 3056.945 52.655 3060.230 54.255 ;
        RECT 3058.360 49.620 3060.230 52.655 ;
        RECT 3028.735 47.805 3032.055 49.405 ;
        RECT 3028.735 47.685 3029.375 47.805 ;
        RECT 2653.830 -3.295 2657.040 -1.770 ;
        RECT 2653.830 -3.370 2657.030 -3.295 ;
      LAYER met5 ;
        RECT 2998.065 4782.790 3001.505 4782.880 ;
        RECT 2998.065 4781.190 3033.895 4782.790 ;
        RECT 2998.065 4781.040 3001.505 4781.190 ;
        RECT 3001.095 4779.260 3004.535 4779.330 ;
        RECT 3030.445 4779.260 3033.885 4779.510 ;
        RECT 3001.095 4777.660 3033.905 4779.260 ;
        RECT 3001.095 4777.490 3004.535 4777.660 ;
        RECT 3004.075 4775.790 3007.515 4775.840 ;
        RECT 3004.075 4774.190 3033.895 4775.790 ;
        RECT 3004.075 4774.000 3007.515 4774.190 ;
        RECT 193.655 4625.595 200.660 4629.595 ;
        RECT 313.655 4625.595 320.660 4629.595 ;
        RECT 433.655 4625.595 440.660 4629.595 ;
        RECT 553.655 4625.595 560.660 4629.595 ;
        RECT 903.655 4625.595 910.660 4629.595 ;
        RECT 1023.655 4625.595 1030.660 4629.595 ;
        RECT 1143.655 4625.595 1150.660 4629.595 ;
        RECT 1263.655 4625.595 1270.660 4629.595 ;
        RECT 1478.655 4625.595 1485.660 4629.595 ;
        RECT 1593.655 4625.595 1600.660 4629.595 ;
        RECT 1958.655 4625.595 1965.660 4629.595 ;
        RECT 2078.655 4625.595 2085.660 4629.595 ;
        RECT 2198.655 4625.595 2205.660 4629.595 ;
        RECT 2318.655 4625.595 2325.660 4629.595 ;
        RECT 2668.655 4625.595 2675.660 4629.595 ;
        RECT 2788.655 4625.595 2795.660 4629.595 ;
        RECT 2908.655 4625.595 2915.660 4629.595 ;
        RECT 2998.095 4625.595 3005.100 4629.595 ;
        RECT -0.815 4514.950 154.345 4516.550 ;
        RECT -0.845 4509.950 152.855 4511.550 ;
        RECT -0.815 4504.950 154.345 4506.550 ;
        RECT 3023.970 4434.840 3179.130 4436.440 ;
        RECT 3025.460 4429.840 3179.160 4431.440 ;
        RECT 3023.970 4424.840 3179.130 4426.440 ;
        RECT -0.815 4409.950 154.345 4411.550 ;
        RECT -0.845 4404.950 152.855 4406.550 ;
        RECT -0.815 4399.950 154.345 4401.550 ;
        RECT 3023.970 4329.850 3179.130 4331.450 ;
        RECT 3025.460 4324.850 3179.160 4326.450 ;
        RECT 3023.970 4319.850 3179.130 4321.450 ;
        RECT -0.815 4304.950 154.345 4306.550 ;
        RECT -0.845 4299.950 152.855 4301.550 ;
        RECT -0.815 4294.950 154.345 4296.550 ;
        RECT 3023.970 4224.850 3179.130 4226.450 ;
        RECT 3025.460 4219.850 3179.160 4221.450 ;
        RECT 3023.970 4214.850 3179.130 4216.450 ;
        RECT -0.815 4199.950 154.345 4201.550 ;
        RECT -0.845 4194.950 152.855 4196.550 ;
        RECT -0.815 4189.950 154.345 4191.550 ;
        RECT 3023.970 4119.850 3179.130 4121.450 ;
        RECT 3025.460 4114.850 3179.160 4116.450 ;
        RECT 3023.970 4109.850 3179.130 4111.450 ;
        RECT 150.450 3996.630 153.890 3996.750 ;
        RECT 1.120 3995.030 153.955 3996.630 ;
        RECT 150.450 3994.910 153.890 3995.030 ;
        RECT 151.755 3991.630 155.195 3991.750 ;
        RECT -1.240 3990.030 155.195 3991.630 ;
        RECT 151.755 3989.910 155.195 3990.030 ;
        RECT 153.015 3986.630 156.455 3986.750 ;
        RECT 1.120 3985.030 156.455 3986.630 ;
        RECT 153.015 3984.910 156.455 3985.030 ;
        RECT 3014.570 3916.065 3018.010 3916.190 ;
        RECT 3014.570 3914.465 3175.305 3916.065 ;
        RECT 3014.570 3914.350 3018.010 3914.465 ;
        RECT 3013.190 3911.065 3016.630 3911.185 ;
        RECT 3013.190 3909.465 3178.610 3911.065 ;
        RECT 3013.190 3909.345 3016.630 3909.465 ;
        RECT 3011.985 3906.065 3015.425 3906.195 ;
        RECT 3011.985 3904.465 3175.305 3906.065 ;
        RECT 3011.985 3904.355 3015.425 3904.465 ;
        RECT 153.010 3891.630 156.450 3891.750 ;
        RECT 1.120 3890.030 156.515 3891.630 ;
        RECT 153.010 3889.910 156.450 3890.030 ;
        RECT 154.320 3886.630 157.760 3886.750 ;
        RECT -1.240 3885.030 157.760 3886.630 ;
        RECT 154.320 3884.910 157.760 3885.030 ;
        RECT 155.575 3881.630 159.015 3881.750 ;
        RECT 1.120 3880.030 159.015 3881.630 ;
        RECT 155.575 3879.910 159.015 3880.030 ;
        RECT 3011.900 3811.065 3015.340 3811.150 ;
        RECT 3011.900 3809.465 3175.305 3811.065 ;
        RECT 3011.900 3809.310 3015.340 3809.465 ;
        RECT 3010.630 3806.065 3014.070 3806.265 ;
        RECT 3010.630 3804.465 3178.610 3806.065 ;
        RECT 3010.630 3804.425 3014.070 3804.465 ;
        RECT 3009.410 3801.065 3012.850 3801.145 ;
        RECT 3009.410 3799.465 3175.305 3801.065 ;
        RECT 3009.410 3799.305 3012.850 3799.465 ;
        RECT 155.575 3786.630 159.015 3786.755 ;
        RECT 1.120 3785.030 159.075 3786.630 ;
        RECT 155.575 3784.915 159.015 3785.030 ;
        RECT 156.875 3781.630 160.315 3781.750 ;
        RECT -1.240 3780.030 160.315 3781.630 ;
        RECT 156.875 3779.910 160.315 3780.030 ;
        RECT 158.130 3776.630 161.570 3776.745 ;
        RECT 1.120 3775.030 161.570 3776.630 ;
        RECT 158.130 3774.905 161.570 3775.030 ;
        RECT 3009.385 3706.065 3012.825 3706.135 ;
        RECT 3009.385 3704.465 3175.305 3706.065 ;
        RECT 3009.385 3704.295 3012.825 3704.465 ;
        RECT 3008.070 3701.065 3011.510 3701.215 ;
        RECT 3008.070 3699.465 3178.610 3701.065 ;
        RECT 3008.070 3699.375 3011.510 3699.465 ;
        RECT 3006.925 3696.065 3010.365 3696.160 ;
        RECT 3006.925 3694.465 3175.305 3696.065 ;
        RECT 3006.925 3694.320 3010.365 3694.465 ;
        RECT 158.135 3681.630 161.575 3681.750 ;
        RECT 1.120 3680.030 161.635 3681.630 ;
        RECT 158.135 3679.910 161.575 3680.030 ;
        RECT 159.440 3676.630 162.880 3676.750 ;
        RECT -1.240 3675.030 162.880 3676.630 ;
        RECT 159.440 3674.910 162.880 3675.030 ;
        RECT 160.700 3671.630 164.140 3671.760 ;
        RECT 1.120 3670.030 164.140 3671.630 ;
        RECT 160.700 3669.920 164.140 3670.030 ;
        RECT 3006.845 3601.065 3010.285 3601.150 ;
        RECT 3006.845 3599.465 3175.305 3601.065 ;
        RECT 3006.845 3599.310 3010.285 3599.465 ;
        RECT 3005.335 3596.065 3008.775 3596.185 ;
        RECT 3005.335 3594.465 3178.605 3596.065 ;
        RECT 3005.335 3594.345 3008.775 3594.465 ;
        RECT 3004.295 3591.065 3007.735 3591.140 ;
        RECT 3004.295 3589.465 3175.305 3591.065 ;
        RECT 3004.295 3589.300 3007.735 3589.465 ;
        RECT 3004.265 3149.955 3007.705 3150.220 ;
        RECT 3004.265 3148.380 3175.305 3149.955 ;
        RECT 3004.615 3148.355 3175.305 3148.380 ;
        RECT 3002.950 3144.955 3006.390 3145.095 ;
        RECT 3002.950 3143.355 3178.605 3144.955 ;
        RECT 3002.950 3143.255 3006.390 3143.355 ;
        RECT 3001.705 3139.955 3005.145 3140.185 ;
        RECT 3001.705 3138.355 3175.305 3139.955 ;
        RECT 3001.705 3138.345 3005.145 3138.355 ;
        RECT 160.695 3027.785 164.135 3027.890 ;
        RECT 1.120 3026.185 164.195 3027.785 ;
        RECT 160.695 3026.050 164.135 3026.185 ;
        RECT 161.995 3022.785 165.435 3022.910 ;
        RECT -1.240 3021.185 165.435 3022.785 ;
        RECT 161.995 3021.070 165.435 3021.185 ;
        RECT 163.260 3017.785 166.700 3017.890 ;
        RECT 1.120 3016.185 166.700 3017.785 ;
        RECT 163.260 3016.050 166.700 3016.185 ;
        RECT 3001.815 2984.955 3005.255 2985.070 ;
        RECT 3001.815 2983.355 3175.305 2984.955 ;
        RECT 3001.815 2983.230 3005.255 2983.355 ;
        RECT 3000.215 2979.955 3003.655 2980.090 ;
        RECT 3000.215 2978.355 3178.605 2979.955 ;
        RECT 3000.215 2978.250 3003.655 2978.355 ;
        RECT 2999.130 2974.955 3002.570 2975.095 ;
        RECT 2999.130 2973.355 3175.305 2974.955 ;
        RECT 2999.130 2973.255 3002.570 2973.355 ;
        RECT 163.260 2862.780 166.700 2862.885 ;
        RECT 1.120 2861.180 166.755 2862.780 ;
        RECT 163.260 2861.045 166.700 2861.180 ;
        RECT 164.555 2857.780 167.995 2857.880 ;
        RECT -1.240 2856.180 167.995 2857.780 ;
        RECT 164.555 2856.040 167.995 2856.180 ;
        RECT 165.815 2852.780 169.255 2852.890 ;
        RECT 1.120 2851.180 169.255 2852.780 ;
        RECT 165.815 2851.050 169.255 2851.180 ;
        RECT 2999.100 2819.955 3002.540 2820.005 ;
        RECT 2999.100 2818.355 3175.305 2819.955 ;
        RECT 2999.100 2818.165 3002.540 2818.355 ;
        RECT 2997.655 2814.955 3001.095 2815.090 ;
        RECT 2997.655 2813.355 3178.605 2814.955 ;
        RECT 2997.655 2813.250 3001.095 2813.355 ;
        RECT 2996.565 2809.955 3000.005 2810.030 ;
        RECT 2996.565 2808.355 3175.305 2809.955 ;
        RECT 2996.565 2808.190 3000.005 2808.355 ;
        RECT 165.820 2697.915 169.260 2698.010 ;
        RECT 1.120 2696.315 169.315 2697.915 ;
        RECT 165.820 2696.170 169.260 2696.315 ;
        RECT 167.115 2692.915 170.555 2693.020 ;
        RECT -0.485 2692.780 170.555 2692.915 ;
        RECT -1.240 2691.315 170.555 2692.780 ;
        RECT -1.240 2691.180 1.565 2691.315 ;
        RECT 167.115 2691.180 170.555 2691.315 ;
        RECT 168.380 2687.915 171.820 2688.025 ;
        RECT 1.120 2686.315 171.820 2687.915 ;
        RECT 168.380 2686.185 171.820 2686.315 ;
        RECT 2996.595 2654.955 3000.035 2655.085 ;
        RECT 2996.595 2653.355 3175.305 2654.955 ;
        RECT 2996.595 2653.245 3000.035 2653.355 ;
        RECT 2995.095 2649.955 2998.535 2650.090 ;
        RECT 2995.095 2648.355 3178.605 2649.955 ;
        RECT 2995.095 2648.250 2998.535 2648.355 ;
        RECT 2994.025 2644.955 2997.465 2645.080 ;
        RECT 2994.025 2643.355 3175.305 2644.955 ;
        RECT 2994.025 2643.240 2997.465 2643.355 ;
        RECT 168.375 2532.780 171.815 2532.885 ;
        RECT 1.120 2531.180 171.875 2532.780 ;
        RECT 168.375 2531.045 171.815 2531.180 ;
        RECT 169.675 2527.780 173.115 2527.895 ;
        RECT -1.240 2526.180 173.115 2527.780 ;
        RECT 169.675 2526.055 173.115 2526.180 ;
        RECT 170.945 2522.780 174.385 2522.890 ;
        RECT 1.120 2521.180 174.385 2522.780 ;
        RECT 170.945 2521.050 174.385 2521.180 ;
        RECT 170.935 2345.665 174.375 2345.790 ;
        RECT 1.120 2344.065 174.435 2345.665 ;
        RECT 170.935 2343.950 174.375 2344.065 ;
        RECT 172.235 2340.665 175.675 2340.785 ;
        RECT -1.240 2339.065 175.675 2340.665 ;
        RECT 172.235 2338.945 175.675 2339.065 ;
        RECT 2994.025 2336.030 2997.465 2336.140 ;
        RECT 173.490 2335.665 176.930 2335.790 ;
        RECT 1.120 2334.065 176.930 2335.665 ;
        RECT 2994.025 2334.430 3175.305 2336.030 ;
        RECT 2994.025 2334.300 2997.465 2334.430 ;
        RECT 173.490 2333.950 176.930 2334.065 ;
        RECT 2992.535 2331.030 2995.975 2331.150 ;
        RECT 2992.535 2329.430 3178.605 2331.030 ;
        RECT 2992.535 2329.310 2995.975 2329.430 ;
        RECT 2991.430 2326.030 2994.870 2326.105 ;
        RECT 2991.430 2324.430 3175.305 2326.030 ;
        RECT 2991.430 2324.265 2994.870 2324.430 ;
        RECT 2991.430 2166.955 2994.870 2167.005 ;
        RECT 2991.430 2165.355 3175.305 2166.955 ;
        RECT 2991.430 2165.165 2994.870 2165.355 ;
        RECT 2989.975 2161.955 2993.415 2162.090 ;
        RECT 2989.975 2160.355 3178.605 2161.955 ;
        RECT 2989.975 2160.250 2993.415 2160.355 ;
        RECT 2988.950 2156.955 2992.390 2157.120 ;
        RECT 2988.950 2155.355 3175.305 2156.955 ;
        RECT 2988.950 2155.280 2992.390 2155.355 ;
        RECT 173.495 2044.780 176.935 2044.885 ;
        RECT 1.120 2043.180 176.995 2044.780 ;
        RECT 173.495 2043.045 176.935 2043.180 ;
        RECT 174.805 2039.780 178.245 2039.895 ;
        RECT -1.240 2038.180 178.245 2039.780 ;
        RECT 174.805 2038.055 178.245 2038.180 ;
        RECT 176.055 2034.780 179.495 2034.895 ;
        RECT 1.120 2033.180 179.495 2034.780 ;
        RECT 176.055 2033.055 179.495 2033.180 ;
        RECT 2988.890 2001.955 2992.330 2002.030 ;
        RECT 2988.890 2000.355 3175.305 2001.955 ;
        RECT 2988.890 2000.190 2992.330 2000.355 ;
        RECT 2987.415 1996.955 2990.855 1997.085 ;
        RECT 2987.415 1995.355 3178.605 1996.955 ;
        RECT 2987.415 1995.245 2990.855 1995.355 ;
        RECT 2986.440 1991.955 2989.880 1992.025 ;
        RECT 2986.440 1990.355 3175.305 1991.955 ;
        RECT 2986.440 1990.185 2989.880 1990.355 ;
        RECT 176.045 1879.780 179.485 1879.880 ;
        RECT 1.120 1878.180 179.555 1879.780 ;
        RECT 176.045 1878.040 179.485 1878.180 ;
        RECT 177.355 1874.780 180.795 1874.880 ;
        RECT -1.240 1873.180 180.795 1874.780 ;
        RECT 177.355 1873.040 180.795 1873.180 ;
        RECT 178.615 1869.780 182.055 1869.880 ;
        RECT 1.120 1868.180 182.055 1869.780 ;
        RECT 178.615 1868.040 182.055 1868.180 ;
        RECT 2986.265 1835.525 2989.705 1835.720 ;
        RECT 2986.265 1833.925 3175.305 1835.525 ;
        RECT 2986.265 1833.880 2989.705 1833.925 ;
        RECT 2984.905 1830.525 2988.345 1830.645 ;
        RECT 3174.725 1830.525 3178.605 1830.670 ;
        RECT 2984.905 1829.070 3178.605 1830.525 ;
        RECT 2984.905 1828.925 3178.445 1829.070 ;
        RECT 2984.905 1828.805 2988.345 1828.925 ;
        RECT 2983.815 1825.525 2987.255 1825.660 ;
        RECT 2983.815 1823.925 3175.305 1825.525 ;
        RECT 2983.815 1823.820 2987.255 1823.925 ;
        RECT 178.615 1716.065 182.055 1716.190 ;
        RECT 1.120 1714.465 182.055 1716.065 ;
        RECT 178.615 1714.350 182.055 1714.465 ;
        RECT 179.915 1711.065 183.355 1711.160 ;
        RECT -1.240 1709.465 183.355 1711.065 ;
        RECT 179.915 1709.320 183.355 1709.465 ;
        RECT 181.180 1706.065 184.620 1706.190 ;
        RECT 1.120 1704.465 184.620 1706.065 ;
        RECT 181.180 1704.350 184.620 1704.465 ;
        RECT 2983.760 1670.670 2987.200 1670.805 ;
        RECT 2983.760 1669.070 3175.305 1670.670 ;
        RECT 2983.760 1668.965 2987.200 1669.070 ;
        RECT 2982.345 1665.670 2985.785 1665.790 ;
        RECT 2982.345 1664.070 3178.605 1665.670 ;
        RECT 2982.345 1663.950 2985.785 1664.070 ;
        RECT 2981.160 1660.670 2984.600 1660.800 ;
        RECT 2981.160 1659.070 3175.305 1660.670 ;
        RECT 2981.160 1658.960 2984.600 1659.070 ;
        RECT 181.055 1551.065 184.495 1551.160 ;
        RECT 1.120 1549.465 184.675 1551.065 ;
        RECT 181.055 1549.320 184.495 1549.465 ;
        RECT 182.475 1546.065 185.915 1546.180 ;
        RECT -1.240 1544.465 185.915 1546.065 ;
        RECT 182.475 1544.340 185.915 1544.465 ;
        RECT 183.655 1541.065 187.095 1541.305 ;
        RECT 1.120 1539.465 187.095 1541.065 ;
        RECT 2641.355 109.285 2644.795 109.410 ;
        RECT 3010.700 109.285 3014.140 109.440 ;
        RECT 2641.355 107.685 3014.140 109.285 ;
        RECT 2641.355 107.570 2644.795 107.685 ;
        RECT 3010.700 107.600 3014.140 107.685 ;
        RECT 2644.710 104.285 2648.150 104.310 ;
        RECT 3011.950 104.285 3015.390 104.395 ;
        RECT 2644.710 102.685 3015.390 104.285 ;
        RECT 2644.710 102.470 2648.150 102.685 ;
        RECT 3011.950 102.555 3015.390 102.685 ;
        RECT 2648.415 99.285 2651.855 99.425 ;
        RECT 3013.180 99.285 3016.620 99.415 ;
        RECT 2648.415 97.685 3016.620 99.285 ;
        RECT 2648.415 97.585 2651.855 97.685 ;
        RECT 3013.180 97.575 3016.620 97.685 ;
        RECT 2651.790 94.285 2655.230 94.350 ;
        RECT 3014.410 94.285 3017.850 94.460 ;
        RECT 2651.790 92.685 3017.850 94.285 ;
        RECT 2651.790 92.510 2655.230 92.685 ;
        RECT 3014.410 92.620 3017.850 92.685 ;
        RECT 2655.445 89.285 2658.885 89.370 ;
        RECT 3015.745 89.285 3019.185 89.395 ;
        RECT 2655.445 87.685 3019.185 89.285 ;
        RECT 2655.445 87.530 2658.885 87.685 ;
        RECT 3015.745 87.555 3019.185 87.685 ;
        RECT 2677.385 84.285 2680.825 84.340 ;
        RECT 3016.995 84.285 3020.435 84.445 ;
        RECT 2677.385 82.685 3020.435 84.285 ;
        RECT 2677.385 82.500 2680.825 82.685 ;
        RECT 3016.995 82.605 3020.435 82.685 ;
        RECT 3018.305 79.285 3021.745 79.480 ;
        RECT 2681.850 77.685 3021.745 79.285 ;
        RECT 3018.305 77.640 3021.745 77.685 ;
        RECT 2679.540 74.285 2682.980 74.370 ;
        RECT 3019.595 74.285 3023.035 74.495 ;
        RECT 2679.540 72.685 3023.035 74.285 ;
        RECT 2679.540 72.530 2682.980 72.685 ;
        RECT 3019.595 72.655 3023.035 72.685 ;
        RECT 3020.800 69.285 3024.240 69.420 ;
        RECT 2683.880 67.685 3024.240 69.285 ;
        RECT 3020.800 67.580 3024.240 67.685 ;
        RECT 2724.440 64.285 2727.880 64.335 ;
        RECT 3022.090 64.285 3025.530 64.455 ;
        RECT 2724.440 62.685 3025.530 64.285 ;
        RECT 2724.440 62.495 2727.880 62.685 ;
        RECT 3022.090 62.615 3025.530 62.685 ;
        RECT 3023.360 59.285 3026.800 59.425 ;
        RECT 2729.310 57.685 3026.800 59.285 ;
        RECT 3023.360 57.585 3026.800 57.685 ;
        RECT 3031.365 59.285 3034.805 59.325 ;
        RECT 3031.365 57.685 3060.265 59.285 ;
        RECT 3031.365 57.485 3034.805 57.685 ;
        RECT 2840.675 54.285 2844.115 54.375 ;
        RECT 3024.740 54.285 3028.180 54.525 ;
        RECT 2840.675 52.685 3028.180 54.285 ;
        RECT 3029.985 54.285 3033.425 54.525 ;
        RECT 3056.825 54.285 3060.265 54.375 ;
        RECT 3029.985 52.685 3060.265 54.285 ;
        RECT 2840.675 52.535 2844.115 52.685 ;
        RECT 3056.825 52.535 3060.265 52.685 ;
        RECT 3028.735 49.285 3032.175 49.525 ;
        RECT 2844.465 47.685 3056.365 49.285 ;
        RECT 2639.760 11.020 2643.200 12.190 ;
        RECT 1451.400 10.350 2643.200 11.020 ;
        RECT 1451.400 9.420 2641.570 10.350 ;
        RECT 2643.185 7.810 2646.625 8.685 ;
        RECT 1451.400 6.845 2646.625 7.810 ;
        RECT 1451.400 6.210 2645.100 6.845 ;
        RECT 2646.695 4.610 2650.135 5.240 ;
        RECT 1451.400 3.400 2650.135 4.610 ;
        RECT 1451.400 3.010 2648.420 3.400 ;
        RECT 2650.120 1.410 2653.560 1.795 ;
        RECT 1451.400 -0.045 2653.560 1.410 ;
        RECT 1451.400 -0.190 2652.500 -0.045 ;
        RECT 2653.710 -1.800 2657.150 -1.650 ;
        RECT 1451.400 -3.400 2657.165 -1.800 ;
        RECT 2653.710 -3.490 2657.150 -3.400 ;
  END
END analog_routes
END LIBRARY

