VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO project_id_rom_32bit
  CLASS BLOCK ;
  FOREIGN project_id_rom_32bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.140 BY 13.680 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 10.135 8.350 10.565 9.135 ;
        RECT 22.555 8.350 22.985 9.135 ;
        RECT 23.015 7.185 23.445 7.970 ;
        RECT 10.135 2.910 10.565 3.695 ;
        RECT 22.555 2.910 22.985 3.695 ;
      LAYER li1 ;
        RECT 0.085 8.995 0.605 9.535 ;
        RECT 26.535 8.995 27.055 9.535 ;
        RECT 0.085 8.245 1.295 8.995 ;
        RECT 2.615 8.245 2.955 8.905 ;
        RECT 3.995 8.245 4.335 8.905 ;
        RECT 5.375 8.245 5.715 8.905 ;
        RECT 6.755 8.245 7.095 8.905 ;
        RECT 8.135 8.245 8.475 8.905 ;
        RECT 9.515 8.245 9.855 8.905 ;
        RECT 10.205 8.245 10.495 8.970 ;
        RECT 11.815 8.245 12.155 8.905 ;
        RECT 13.195 8.245 13.535 8.905 ;
        RECT 14.575 8.245 14.915 8.905 ;
        RECT 16.415 8.245 16.755 8.905 ;
        RECT 17.795 8.245 18.135 8.905 ;
        RECT 19.175 8.245 19.515 8.905 ;
        RECT 20.555 8.245 20.895 8.905 ;
        RECT 21.935 8.245 22.275 8.905 ;
        RECT 22.625 8.245 22.915 8.970 ;
        RECT 23.775 8.245 24.115 8.905 ;
        RECT 25.155 8.245 25.495 8.905 ;
        RECT 25.845 8.245 27.055 8.995 ;
        RECT 0.000 8.075 27.140 8.245 ;
        RECT 0.085 7.325 1.295 8.075 ;
        RECT 0.085 6.785 0.605 7.325 ;
        RECT 1.465 7.305 4.055 8.075 ;
        RECT 4.225 7.305 9.570 8.075 ;
        RECT 9.745 7.305 15.090 8.075 ;
        RECT 15.265 7.305 20.610 8.075 ;
        RECT 20.785 7.305 22.455 8.075 ;
        RECT 23.085 7.350 23.375 8.075 ;
        RECT 23.545 7.305 25.215 8.075 ;
        RECT 25.845 7.325 27.055 8.075 ;
        RECT 1.465 6.785 2.675 7.305 ;
        RECT 4.225 6.785 6.805 7.305 ;
        RECT 9.745 6.785 12.325 7.305 ;
        RECT 15.265 6.785 17.845 7.305 ;
        RECT 20.785 6.785 21.535 7.305 ;
        RECT 23.545 6.785 24.295 7.305 ;
        RECT 26.535 6.785 27.055 7.325 ;
        RECT 0.085 3.555 0.605 4.095 ;
        RECT 26.535 3.555 27.055 4.095 ;
        RECT 0.085 2.805 1.295 3.555 ;
        RECT 2.615 2.805 2.955 3.465 ;
        RECT 3.995 2.805 4.335 3.465 ;
        RECT 5.375 2.805 5.715 3.465 ;
        RECT 6.755 2.805 7.095 3.465 ;
        RECT 8.135 2.805 8.475 3.465 ;
        RECT 9.515 2.805 9.855 3.465 ;
        RECT 10.205 2.805 10.495 3.530 ;
        RECT 11.815 2.805 12.155 3.465 ;
        RECT 13.195 2.805 13.535 3.465 ;
        RECT 14.575 2.805 14.915 3.465 ;
        RECT 16.415 2.805 16.755 3.465 ;
        RECT 17.795 2.805 18.135 3.465 ;
        RECT 19.175 2.805 19.515 3.465 ;
        RECT 20.555 2.805 20.895 3.465 ;
        RECT 21.935 2.805 22.275 3.465 ;
        RECT 22.625 2.805 22.915 3.530 ;
        RECT 23.775 2.805 24.115 3.465 ;
        RECT 25.155 2.805 25.495 3.465 ;
        RECT 25.845 2.805 27.055 3.555 ;
        RECT 0.000 2.635 27.140 2.805 ;
      LAYER met1 ;
        RECT 0.000 7.920 27.140 8.400 ;
        RECT 0.000 2.480 27.140 2.960 ;
      LAYER met2 ;
        RECT 1.130 7.920 2.350 8.400 ;
        RECT 8.130 7.920 9.350 8.400 ;
        RECT 15.130 7.920 16.350 8.400 ;
        RECT 22.130 7.920 23.350 8.400 ;
        RECT 1.290 2.960 1.830 7.920 ;
        RECT 1.130 2.480 2.350 2.960 ;
        RECT 8.130 2.480 9.350 2.960 ;
        RECT 15.130 2.480 16.350 2.960 ;
        RECT 22.130 2.480 23.350 2.960 ;
      LAYER met3 ;
        RECT 1.040 7.920 23.440 8.400 ;
        RECT 1.040 2.480 23.440 2.960 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 9.465 27.330 11.070 ;
        RECT -0.190 4.025 27.330 6.855 ;
      LAYER li1 ;
        RECT 0.000 10.795 27.140 10.965 ;
        RECT 0.085 9.705 1.295 10.795 ;
        RECT 2.115 10.070 2.445 10.795 ;
        RECT 3.495 10.070 3.825 10.795 ;
        RECT 4.875 10.070 5.205 10.795 ;
        RECT 6.255 10.070 6.585 10.795 ;
        RECT 7.635 10.070 7.965 10.795 ;
        RECT 9.015 10.070 9.345 10.795 ;
        RECT 0.775 9.165 1.295 9.705 ;
        RECT 10.205 9.630 10.495 10.795 ;
        RECT 11.315 10.070 11.645 10.795 ;
        RECT 12.695 10.070 13.025 10.795 ;
        RECT 14.075 10.070 14.405 10.795 ;
        RECT 15.915 10.070 16.245 10.795 ;
        RECT 17.295 10.070 17.625 10.795 ;
        RECT 18.675 10.070 19.005 10.795 ;
        RECT 20.055 10.070 20.385 10.795 ;
        RECT 21.435 10.070 21.765 10.795 ;
        RECT 22.625 9.630 22.915 10.795 ;
        RECT 23.275 10.070 23.605 10.795 ;
        RECT 24.655 10.070 24.985 10.795 ;
        RECT 25.845 9.705 27.055 10.795 ;
        RECT 25.845 9.165 26.365 9.705 ;
        RECT 0.775 6.615 1.295 7.155 ;
        RECT 2.845 6.615 4.055 7.135 ;
        RECT 6.975 6.615 9.570 7.135 ;
        RECT 12.495 6.615 15.090 7.135 ;
        RECT 18.015 6.615 20.610 7.135 ;
        RECT 21.705 6.615 22.455 7.135 ;
        RECT 0.085 5.525 1.295 6.615 ;
        RECT 1.465 5.525 4.055 6.615 ;
        RECT 4.225 5.525 9.570 6.615 ;
        RECT 9.745 5.525 15.090 6.615 ;
        RECT 15.265 5.525 20.610 6.615 ;
        RECT 20.785 5.525 22.455 6.615 ;
        RECT 23.085 5.525 23.375 6.690 ;
        RECT 24.465 6.615 25.215 7.135 ;
        RECT 23.545 5.525 25.215 6.615 ;
        RECT 25.845 6.615 26.365 7.155 ;
        RECT 25.845 5.525 27.055 6.615 ;
        RECT 0.000 5.355 27.140 5.525 ;
        RECT 0.085 4.265 1.295 5.355 ;
        RECT 2.115 4.630 2.445 5.355 ;
        RECT 3.495 4.630 3.825 5.355 ;
        RECT 4.875 4.630 5.205 5.355 ;
        RECT 6.255 4.630 6.585 5.355 ;
        RECT 7.635 4.630 7.965 5.355 ;
        RECT 9.015 4.630 9.345 5.355 ;
        RECT 0.775 3.725 1.295 4.265 ;
        RECT 10.205 4.190 10.495 5.355 ;
        RECT 11.315 4.630 11.645 5.355 ;
        RECT 12.695 4.630 13.025 5.355 ;
        RECT 14.075 4.630 14.405 5.355 ;
        RECT 15.915 4.630 16.245 5.355 ;
        RECT 17.295 4.630 17.625 5.355 ;
        RECT 18.675 4.630 19.005 5.355 ;
        RECT 20.055 4.630 20.385 5.355 ;
        RECT 21.435 4.630 21.765 5.355 ;
        RECT 22.625 4.190 22.915 5.355 ;
        RECT 23.275 4.630 23.605 5.355 ;
        RECT 24.655 4.630 24.985 5.355 ;
        RECT 25.845 4.265 27.055 5.355 ;
        RECT 25.845 3.725 26.365 4.265 ;
      LAYER met1 ;
        RECT 0.000 10.640 27.140 11.120 ;
        RECT 0.000 5.200 27.140 5.680 ;
      LAYER met2 ;
        RECT 4.630 10.640 5.850 11.120 ;
        RECT 11.630 10.640 12.850 11.120 ;
        RECT 18.630 10.640 19.850 11.120 ;
        RECT 4.790 5.680 5.330 10.640 ;
        RECT 4.630 5.200 5.850 5.680 ;
        RECT 11.630 5.200 12.850 5.680 ;
        RECT 18.630 5.200 19.850 5.680 ;
      LAYER met3 ;
        RECT 4.540 10.640 19.940 11.120 ;
        RECT 4.540 5.200 19.940 5.680 ;
    END
  END VPWR
  PIN gpio_defaults[0]
    PORT
      LAYER li1 ;
        RECT 2.615 3.635 3.135 5.185 ;
      LAYER met1 ;
        RECT 2.035 3.980 2.325 4.025 ;
        RECT 2.725 3.980 3.015 4.025 ;
        RECT 2.035 3.840 3.015 3.980 ;
        RECT 2.035 3.795 2.325 3.840 ;
        RECT 2.725 3.795 3.015 3.840 ;
        RECT 2.815 3.555 2.955 3.795 ;
        RECT 2.770 3.235 3.030 3.555 ;
      LAYER met2 ;
        RECT 2.740 3.465 3.060 3.525 ;
        RECT 2.610 3.265 3.060 3.465 ;
        RECT 2.610 2.370 2.750 3.265 ;
        RECT 2.455 2.225 2.750 2.370 ;
        RECT 2.455 2.000 2.595 2.225 ;
        RECT 2.390 0.000 2.670 2.000 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[1]
    PORT
      LAYER li1 ;
        RECT 2.615 9.075 3.135 10.625 ;
      LAYER met1 ;
        RECT 2.770 9.785 3.030 10.105 ;
        RECT 2.815 9.545 2.955 9.785 ;
        RECT 2.035 9.500 2.325 9.545 ;
        RECT 2.725 9.500 3.015 9.545 ;
        RECT 2.035 9.360 3.015 9.500 ;
        RECT 2.035 9.315 2.325 9.360 ;
        RECT 2.725 9.315 3.015 9.360 ;
      LAYER met2 ;
        RECT 2.390 11.680 2.670 13.680 ;
        RECT 2.450 10.015 2.590 11.680 ;
        RECT 2.735 10.015 3.060 10.075 ;
        RECT 2.450 9.875 3.060 10.015 ;
        RECT 2.735 9.815 3.060 9.875 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[2]
    PORT
      LAYER li1 ;
        RECT 3.995 3.635 4.515 5.185 ;
      LAYER met1 ;
        RECT 3.415 3.980 3.705 4.025 ;
        RECT 4.105 3.980 4.395 4.025 ;
        RECT 3.415 3.840 4.395 3.980 ;
        RECT 3.415 3.795 3.705 3.840 ;
        RECT 4.105 3.795 4.395 3.840 ;
        RECT 4.195 3.555 4.335 3.795 ;
        RECT 4.150 3.235 4.410 3.555 ;
      LAYER met2 ;
        RECT 4.120 3.465 4.440 3.525 ;
        RECT 3.840 3.325 4.440 3.465 ;
        RECT 3.840 2.000 3.980 3.325 ;
        RECT 4.120 3.265 4.440 3.325 ;
        RECT 3.770 0.000 4.050 2.000 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[3]
    PORT
      LAYER li1 ;
        RECT 3.995 9.075 4.515 10.625 ;
      LAYER met1 ;
        RECT 4.150 9.785 4.410 10.105 ;
        RECT 4.195 9.545 4.335 9.785 ;
        RECT 3.415 9.500 3.705 9.545 ;
        RECT 4.105 9.500 4.395 9.545 ;
        RECT 3.415 9.360 4.395 9.500 ;
        RECT 3.415 9.315 3.705 9.360 ;
        RECT 4.105 9.315 4.395 9.360 ;
      LAYER met2 ;
        RECT 3.770 11.680 4.050 13.680 ;
        RECT 3.840 10.015 3.980 11.680 ;
        RECT 4.120 10.015 4.440 10.075 ;
        RECT 3.840 9.875 4.440 10.015 ;
        RECT 4.120 9.815 4.440 9.875 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[4]
    PORT
      LAYER li1 ;
        RECT 5.375 3.635 5.895 5.185 ;
      LAYER met1 ;
        RECT 4.795 3.980 5.085 4.025 ;
        RECT 5.485 3.980 5.775 4.025 ;
        RECT 4.795 3.840 5.775 3.980 ;
        RECT 4.795 3.795 5.085 3.840 ;
        RECT 5.485 3.795 5.775 3.840 ;
        RECT 5.575 3.555 5.715 3.795 ;
        RECT 5.530 3.235 5.790 3.555 ;
      LAYER met2 ;
        RECT 5.500 3.465 5.820 3.525 ;
        RECT 5.220 3.325 5.820 3.465 ;
        RECT 5.220 2.000 5.360 3.325 ;
        RECT 5.500 3.265 5.820 3.325 ;
        RECT 5.150 0.000 5.430 2.000 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[5]
    PORT
      LAYER li1 ;
        RECT 5.375 9.075 5.895 10.625 ;
      LAYER met1 ;
        RECT 5.530 9.785 5.790 10.105 ;
        RECT 5.575 9.545 5.715 9.785 ;
        RECT 4.795 9.500 5.085 9.545 ;
        RECT 5.485 9.500 5.775 9.545 ;
        RECT 4.795 9.360 5.775 9.500 ;
        RECT 4.795 9.315 5.085 9.360 ;
        RECT 5.485 9.315 5.775 9.360 ;
      LAYER met2 ;
        RECT 5.150 11.680 5.430 13.680 ;
        RECT 5.215 11.505 5.355 11.680 ;
        RECT 5.215 11.365 6.190 11.505 ;
        RECT 5.500 10.015 5.820 10.075 ;
        RECT 6.050 10.015 6.190 11.365 ;
        RECT 5.500 9.875 6.190 10.015 ;
        RECT 5.500 9.815 5.820 9.875 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[6]
    PORT
      LAYER li1 ;
        RECT 6.755 3.635 7.275 5.185 ;
      LAYER met1 ;
        RECT 6.175 3.980 6.465 4.025 ;
        RECT 6.865 3.980 7.155 4.025 ;
        RECT 6.175 3.840 7.155 3.980 ;
        RECT 6.175 3.795 6.465 3.840 ;
        RECT 6.865 3.795 7.155 3.840 ;
        RECT 6.955 3.555 7.095 3.795 ;
        RECT 6.910 3.235 7.170 3.555 ;
      LAYER met2 ;
        RECT 6.880 3.465 7.200 3.525 ;
        RECT 6.600 3.325 7.200 3.465 ;
        RECT 6.600 2.000 6.740 3.325 ;
        RECT 6.880 3.265 7.200 3.325 ;
        RECT 6.530 0.000 6.810 2.000 ;
    END
  END gpio_defaults[6]
  PIN gpio_defaults[7]
    PORT
      LAYER li1 ;
        RECT 6.755 9.075 7.275 10.625 ;
      LAYER met1 ;
        RECT 6.910 9.785 7.170 10.105 ;
        RECT 6.955 9.545 7.095 9.785 ;
        RECT 6.175 9.500 6.465 9.545 ;
        RECT 6.865 9.500 7.155 9.545 ;
        RECT 6.175 9.360 7.155 9.500 ;
        RECT 6.175 9.315 6.465 9.360 ;
        RECT 6.865 9.315 7.155 9.360 ;
      LAYER met2 ;
        RECT 6.530 11.680 6.810 13.680 ;
        RECT 6.600 10.015 6.740 11.680 ;
        RECT 6.880 10.015 7.200 10.075 ;
        RECT 6.600 9.875 7.200 10.015 ;
        RECT 6.880 9.815 7.200 9.875 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[8]
    PORT
      LAYER li1 ;
        RECT 8.135 3.635 8.655 5.185 ;
      LAYER met1 ;
        RECT 7.555 3.980 7.845 4.025 ;
        RECT 8.245 3.980 8.535 4.025 ;
        RECT 7.555 3.840 8.535 3.980 ;
        RECT 7.555 3.795 7.845 3.840 ;
        RECT 8.245 3.795 8.535 3.840 ;
        RECT 8.335 3.555 8.475 3.795 ;
        RECT 8.290 3.235 8.550 3.555 ;
      LAYER met2 ;
        RECT 8.260 3.465 8.580 3.525 ;
        RECT 7.780 3.325 8.580 3.465 ;
        RECT 7.780 2.325 7.920 3.325 ;
        RECT 8.260 3.265 8.580 3.325 ;
        RECT 7.780 2.185 8.120 2.325 ;
        RECT 7.980 2.000 8.120 2.185 ;
        RECT 7.910 0.000 8.190 2.000 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[9]
    PORT
      LAYER li1 ;
        RECT 8.135 9.075 8.655 10.625 ;
      LAYER met1 ;
        RECT 8.290 9.785 8.550 10.105 ;
        RECT 8.335 9.545 8.475 9.785 ;
        RECT 7.555 9.500 7.845 9.545 ;
        RECT 8.245 9.500 8.535 9.545 ;
        RECT 7.555 9.360 8.535 9.500 ;
        RECT 7.555 9.315 7.845 9.360 ;
        RECT 8.245 9.315 8.535 9.360 ;
      LAYER met2 ;
        RECT 7.910 11.680 8.190 13.680 ;
        RECT 7.965 10.015 8.105 11.680 ;
        RECT 8.260 10.015 8.580 10.075 ;
        RECT 7.965 9.875 8.580 10.015 ;
        RECT 8.260 9.815 8.580 9.875 ;
    END
  END gpio_defaults[9]
  PIN gpio_defaults[10]
    PORT
      LAYER li1 ;
        RECT 9.515 3.635 10.035 5.185 ;
      LAYER met1 ;
        RECT 8.935 3.980 9.225 4.025 ;
        RECT 9.625 3.980 9.915 4.025 ;
        RECT 8.935 3.840 9.915 3.980 ;
        RECT 8.935 3.795 9.225 3.840 ;
        RECT 9.625 3.795 9.915 3.840 ;
        RECT 9.715 3.555 9.855 3.795 ;
        RECT 9.670 3.235 9.930 3.555 ;
      LAYER met2 ;
        RECT 9.640 3.265 9.960 3.525 ;
        RECT 9.725 2.415 9.865 3.265 ;
        RECT 9.725 2.265 9.960 2.415 ;
        RECT 9.820 2.000 9.960 2.265 ;
        RECT 9.750 0.000 10.030 2.000 ;
    END
  END gpio_defaults[10]
  PIN gpio_defaults[11]
    PORT
      LAYER li1 ;
        RECT 9.515 9.075 10.035 10.625 ;
      LAYER met1 ;
        RECT 9.670 9.785 9.930 10.105 ;
        RECT 9.715 9.545 9.855 9.785 ;
        RECT 8.935 9.500 9.225 9.545 ;
        RECT 9.625 9.500 9.915 9.545 ;
        RECT 8.935 9.360 9.915 9.500 ;
        RECT 8.935 9.315 9.225 9.360 ;
        RECT 9.625 9.315 9.915 9.360 ;
      LAYER met2 ;
        RECT 9.750 11.680 10.030 13.680 ;
        RECT 9.815 11.260 9.955 11.680 ;
        RECT 9.725 11.120 9.955 11.260 ;
        RECT 9.725 10.075 9.865 11.120 ;
        RECT 9.640 9.815 9.960 10.075 ;
    END
  END gpio_defaults[11]
  PIN gpio_defaults[12]
    PORT
      LAYER li1 ;
        RECT 11.815 3.635 12.335 5.185 ;
      LAYER met1 ;
        RECT 11.235 3.980 11.525 4.025 ;
        RECT 11.925 3.980 12.215 4.025 ;
        RECT 11.235 3.840 12.215 3.980 ;
        RECT 11.235 3.795 11.525 3.840 ;
        RECT 11.925 3.795 12.215 3.840 ;
        RECT 12.015 3.555 12.155 3.795 ;
        RECT 11.970 3.235 12.230 3.555 ;
      LAYER met2 ;
        RECT 11.940 3.465 12.260 3.525 ;
        RECT 11.660 3.325 12.260 3.465 ;
        RECT 11.660 2.000 11.800 3.325 ;
        RECT 11.940 3.265 12.260 3.325 ;
        RECT 11.590 0.000 11.870 2.000 ;
    END
  END gpio_defaults[12]
  PIN gpio_defaults[13]
    PORT
      LAYER li1 ;
        RECT 11.815 9.075 12.335 10.625 ;
      LAYER met1 ;
        RECT 11.970 9.785 12.230 10.105 ;
        RECT 12.015 9.545 12.155 9.785 ;
        RECT 11.235 9.500 11.525 9.545 ;
        RECT 11.925 9.500 12.215 9.545 ;
        RECT 11.235 9.360 12.215 9.500 ;
        RECT 11.235 9.315 11.525 9.360 ;
        RECT 11.925 9.315 12.215 9.360 ;
      LAYER met2 ;
        RECT 11.590 11.680 11.870 13.680 ;
        RECT 11.650 11.485 11.790 11.680 ;
        RECT 11.250 11.345 11.790 11.485 ;
        RECT 11.250 10.015 11.390 11.345 ;
        RECT 11.940 10.015 12.260 10.075 ;
        RECT 11.250 9.875 12.260 10.015 ;
        RECT 11.940 9.815 12.260 9.875 ;
    END
  END gpio_defaults[13]
  PIN gpio_defaults[14]
    PORT
      LAYER li1 ;
        RECT 13.195 3.635 13.715 5.185 ;
      LAYER met1 ;
        RECT 12.615 3.980 12.905 4.025 ;
        RECT 13.305 3.980 13.595 4.025 ;
        RECT 12.615 3.840 13.595 3.980 ;
        RECT 12.615 3.795 12.905 3.840 ;
        RECT 13.305 3.795 13.595 3.840 ;
        RECT 13.395 3.555 13.535 3.795 ;
        RECT 13.350 3.235 13.610 3.555 ;
      LAYER met2 ;
        RECT 13.320 3.465 13.640 3.525 ;
        RECT 13.040 3.325 13.640 3.465 ;
        RECT 13.040 2.000 13.180 3.325 ;
        RECT 13.320 3.265 13.640 3.325 ;
        RECT 12.970 0.000 13.250 2.000 ;
    END
  END gpio_defaults[14]
  PIN gpio_defaults[15]
    PORT
      LAYER li1 ;
        RECT 13.195 9.075 13.715 10.625 ;
      LAYER met1 ;
        RECT 13.350 9.785 13.610 10.105 ;
        RECT 13.395 9.545 13.535 9.785 ;
        RECT 12.615 9.500 12.905 9.545 ;
        RECT 13.305 9.500 13.595 9.545 ;
        RECT 12.615 9.360 13.595 9.500 ;
        RECT 12.615 9.315 12.905 9.360 ;
        RECT 13.305 9.315 13.595 9.360 ;
      LAYER met2 ;
        RECT 12.970 11.680 13.250 13.680 ;
        RECT 13.040 10.015 13.180 11.680 ;
        RECT 13.320 10.015 13.640 10.075 ;
        RECT 13.040 9.875 13.640 10.015 ;
        RECT 13.320 9.815 13.640 9.875 ;
    END
  END gpio_defaults[15]
  PIN gpio_defaults[16]
    PORT
      LAYER li1 ;
        RECT 14.575 3.635 15.095 5.185 ;
      LAYER met1 ;
        RECT 13.995 3.980 14.285 4.025 ;
        RECT 14.685 3.980 14.975 4.025 ;
        RECT 13.995 3.840 14.975 3.980 ;
        RECT 13.995 3.795 14.285 3.840 ;
        RECT 14.685 3.795 14.975 3.840 ;
        RECT 14.775 3.555 14.915 3.795 ;
        RECT 14.730 3.235 14.990 3.555 ;
      LAYER met2 ;
        RECT 14.700 3.465 15.020 3.525 ;
        RECT 14.420 3.325 15.020 3.465 ;
        RECT 14.420 2.000 14.560 3.325 ;
        RECT 14.700 3.265 15.020 3.325 ;
        RECT 14.350 0.000 14.630 2.000 ;
    END
  END gpio_defaults[16]
  PIN gpio_defaults[17]
    PORT
      LAYER li1 ;
        RECT 14.575 9.075 15.095 10.625 ;
      LAYER met1 ;
        RECT 14.730 9.785 14.990 10.105 ;
        RECT 14.775 9.545 14.915 9.785 ;
        RECT 13.995 9.500 14.285 9.545 ;
        RECT 14.685 9.500 14.975 9.545 ;
        RECT 13.995 9.360 14.975 9.500 ;
        RECT 13.995 9.315 14.285 9.360 ;
        RECT 14.685 9.315 14.975 9.360 ;
      LAYER met2 ;
        RECT 14.350 11.680 14.630 13.680 ;
        RECT 14.420 10.015 14.560 11.680 ;
        RECT 14.700 10.015 15.020 10.075 ;
        RECT 14.420 9.875 15.020 10.015 ;
        RECT 14.700 9.815 15.020 9.875 ;
    END
  END gpio_defaults[17]
  PIN gpio_defaults[18]
    PORT
      LAYER li1 ;
        RECT 16.415 3.635 16.935 5.185 ;
      LAYER met1 ;
        RECT 15.835 3.980 16.125 4.025 ;
        RECT 16.525 3.980 16.815 4.025 ;
        RECT 15.835 3.840 16.815 3.980 ;
        RECT 15.835 3.795 16.125 3.840 ;
        RECT 16.525 3.795 16.815 3.840 ;
        RECT 16.595 3.555 16.735 3.795 ;
        RECT 16.550 3.235 16.810 3.555 ;
      LAYER met2 ;
        RECT 16.520 3.265 16.840 3.525 ;
        RECT 16.600 2.295 16.740 3.265 ;
        RECT 16.260 2.155 16.740 2.295 ;
        RECT 16.260 2.000 16.400 2.155 ;
        RECT 16.190 0.000 16.470 2.000 ;
    END
  END gpio_defaults[18]
  PIN gpio_defaults[19]
    PORT
      LAYER li1 ;
        RECT 16.415 9.075 16.935 10.625 ;
      LAYER met1 ;
        RECT 16.550 9.785 16.810 10.105 ;
        RECT 16.595 9.545 16.735 9.785 ;
        RECT 15.835 9.500 16.125 9.545 ;
        RECT 16.525 9.500 16.815 9.545 ;
        RECT 15.835 9.360 16.815 9.500 ;
        RECT 15.835 9.315 16.125 9.360 ;
        RECT 16.525 9.315 16.815 9.360 ;
      LAYER met2 ;
        RECT 16.190 11.680 16.470 13.680 ;
        RECT 16.245 10.370 16.385 11.680 ;
        RECT 16.245 10.230 16.740 10.370 ;
        RECT 16.600 10.075 16.740 10.230 ;
        RECT 16.520 9.815 16.840 10.075 ;
    END
  END gpio_defaults[19]
  PIN gpio_defaults[20]
    PORT
      LAYER li1 ;
        RECT 17.795 3.635 18.315 5.185 ;
      LAYER met1 ;
        RECT 17.215 3.980 17.505 4.025 ;
        RECT 17.905 3.980 18.195 4.025 ;
        RECT 17.215 3.840 18.195 3.980 ;
        RECT 17.215 3.795 17.505 3.840 ;
        RECT 17.905 3.795 18.195 3.840 ;
        RECT 17.995 3.555 18.135 3.795 ;
        RECT 17.950 3.235 18.210 3.555 ;
      LAYER met2 ;
        RECT 17.920 3.465 18.240 3.525 ;
        RECT 17.640 3.325 18.240 3.465 ;
        RECT 17.640 2.000 17.780 3.325 ;
        RECT 17.920 3.265 18.240 3.325 ;
        RECT 17.570 0.000 17.850 2.000 ;
    END
  END gpio_defaults[20]
  PIN gpio_defaults[21]
    PORT
      LAYER li1 ;
        RECT 17.795 9.075 18.315 10.625 ;
      LAYER met1 ;
        RECT 17.950 9.785 18.210 10.105 ;
        RECT 17.995 9.545 18.135 9.785 ;
        RECT 17.215 9.500 17.505 9.545 ;
        RECT 17.905 9.500 18.195 9.545 ;
        RECT 17.215 9.360 18.195 9.500 ;
        RECT 17.215 9.315 17.505 9.360 ;
        RECT 17.905 9.315 18.195 9.360 ;
      LAYER met2 ;
        RECT 17.570 11.680 17.850 13.680 ;
        RECT 17.640 10.015 17.780 11.680 ;
        RECT 17.920 10.015 18.240 10.075 ;
        RECT 17.640 9.875 18.240 10.015 ;
        RECT 17.920 9.815 18.240 9.875 ;
    END
  END gpio_defaults[21]
  PIN gpio_defaults[22]
    PORT
      LAYER li1 ;
        RECT 19.175 3.635 19.695 5.185 ;
      LAYER met1 ;
        RECT 18.595 3.980 18.885 4.025 ;
        RECT 19.285 3.980 19.575 4.025 ;
        RECT 18.595 3.840 19.575 3.980 ;
        RECT 18.595 3.795 18.885 3.840 ;
        RECT 19.285 3.795 19.575 3.840 ;
        RECT 19.375 3.555 19.515 3.795 ;
        RECT 19.330 3.235 19.590 3.555 ;
      LAYER met2 ;
        RECT 19.300 3.465 19.620 3.525 ;
        RECT 19.020 3.325 19.620 3.465 ;
        RECT 19.020 2.000 19.160 3.325 ;
        RECT 19.300 3.265 19.620 3.325 ;
        RECT 18.950 0.000 19.230 2.000 ;
    END
  END gpio_defaults[22]
  PIN gpio_defaults[23]
    PORT
      LAYER li1 ;
        RECT 19.175 9.075 19.695 10.625 ;
      LAYER met1 ;
        RECT 19.330 9.785 19.590 10.105 ;
        RECT 19.375 9.545 19.515 9.785 ;
        RECT 18.595 9.500 18.885 9.545 ;
        RECT 19.285 9.500 19.575 9.545 ;
        RECT 18.595 9.360 19.575 9.500 ;
        RECT 18.595 9.315 18.885 9.360 ;
        RECT 19.285 9.315 19.575 9.360 ;
      LAYER met2 ;
        RECT 18.950 11.680 19.230 13.680 ;
        RECT 19.015 11.495 19.155 11.680 ;
        RECT 19.015 11.355 20.175 11.495 ;
        RECT 19.300 10.015 19.620 10.075 ;
        RECT 20.035 10.015 20.175 11.355 ;
        RECT 19.300 9.875 20.175 10.015 ;
        RECT 19.300 9.815 19.620 9.875 ;
    END
  END gpio_defaults[23]
  PIN gpio_defaults[24]
    PORT
      LAYER li1 ;
        RECT 20.555 3.635 21.075 5.185 ;
      LAYER met1 ;
        RECT 19.975 3.980 20.265 4.025 ;
        RECT 20.665 3.980 20.955 4.025 ;
        RECT 19.975 3.840 20.955 3.980 ;
        RECT 19.975 3.795 20.265 3.840 ;
        RECT 20.665 3.795 20.955 3.840 ;
        RECT 20.755 3.555 20.895 3.795 ;
        RECT 20.710 3.235 20.970 3.555 ;
      LAYER met2 ;
        RECT 20.680 3.465 21.000 3.525 ;
        RECT 20.400 3.325 21.000 3.465 ;
        RECT 20.400 2.000 20.540 3.325 ;
        RECT 20.680 3.265 21.000 3.325 ;
        RECT 20.330 0.000 20.610 2.000 ;
    END
  END gpio_defaults[24]
  PIN gpio_defaults[25]
    PORT
      LAYER li1 ;
        RECT 20.555 9.075 21.075 10.625 ;
      LAYER met1 ;
        RECT 20.710 9.785 20.970 10.105 ;
        RECT 20.755 9.545 20.895 9.785 ;
        RECT 19.975 9.500 20.265 9.545 ;
        RECT 20.665 9.500 20.955 9.545 ;
        RECT 19.975 9.360 20.955 9.500 ;
        RECT 19.975 9.315 20.265 9.360 ;
        RECT 20.665 9.315 20.955 9.360 ;
      LAYER met2 ;
        RECT 20.330 11.680 20.610 13.680 ;
        RECT 20.400 10.015 20.540 11.680 ;
        RECT 20.680 10.015 21.000 10.075 ;
        RECT 20.400 9.875 21.000 10.015 ;
        RECT 20.680 9.815 21.000 9.875 ;
    END
  END gpio_defaults[25]
  PIN gpio_defaults[26]
    PORT
      LAYER li1 ;
        RECT 21.935 3.635 22.455 5.185 ;
      LAYER met1 ;
        RECT 21.355 3.980 21.645 4.025 ;
        RECT 22.045 3.980 22.335 4.025 ;
        RECT 21.355 3.840 22.335 3.980 ;
        RECT 21.355 3.795 21.645 3.840 ;
        RECT 22.045 3.795 22.335 3.840 ;
        RECT 22.135 3.555 22.275 3.795 ;
        RECT 22.090 3.235 22.350 3.555 ;
      LAYER met2 ;
        RECT 22.060 3.465 22.380 3.525 ;
        RECT 21.780 3.325 22.380 3.465 ;
        RECT 21.780 2.000 21.920 3.325 ;
        RECT 22.060 3.265 22.380 3.325 ;
        RECT 21.710 0.000 21.990 2.000 ;
    END
  END gpio_defaults[26]
  PIN gpio_defaults[27]
    PORT
      LAYER li1 ;
        RECT 21.935 9.075 22.455 10.625 ;
      LAYER met1 ;
        RECT 22.090 9.785 22.350 10.105 ;
        RECT 22.135 9.545 22.275 9.785 ;
        RECT 21.355 9.500 21.645 9.545 ;
        RECT 22.045 9.500 22.335 9.545 ;
        RECT 21.355 9.360 22.335 9.500 ;
        RECT 21.355 9.315 21.645 9.360 ;
        RECT 22.045 9.315 22.335 9.360 ;
      LAYER met2 ;
        RECT 21.710 11.680 21.990 13.680 ;
        RECT 21.780 10.015 21.920 11.680 ;
        RECT 22.060 10.015 22.380 10.075 ;
        RECT 21.780 9.875 22.380 10.015 ;
        RECT 22.060 9.815 22.380 9.875 ;
    END
  END gpio_defaults[27]
  PIN gpio_defaults[28]
    PORT
      LAYER li1 ;
        RECT 23.775 3.635 24.295 5.185 ;
      LAYER met1 ;
        RECT 23.195 3.980 23.485 4.025 ;
        RECT 23.885 3.980 24.175 4.025 ;
        RECT 23.195 3.840 24.175 3.980 ;
        RECT 23.195 3.795 23.485 3.840 ;
        RECT 23.885 3.795 24.175 3.840 ;
        RECT 23.975 3.555 24.115 3.795 ;
        RECT 23.930 3.235 24.190 3.555 ;
      LAYER met2 ;
        RECT 23.900 3.465 24.220 3.525 ;
        RECT 23.620 3.325 24.220 3.465 ;
        RECT 23.620 2.000 23.760 3.325 ;
        RECT 23.900 3.265 24.220 3.325 ;
        RECT 23.550 0.000 23.830 2.000 ;
    END
  END gpio_defaults[28]
  PIN gpio_defaults[29]
    PORT
      LAYER li1 ;
        RECT 23.775 9.075 24.295 10.625 ;
      LAYER met1 ;
        RECT 23.930 9.785 24.190 10.105 ;
        RECT 23.975 9.545 24.115 9.785 ;
        RECT 23.195 9.500 23.485 9.545 ;
        RECT 23.885 9.500 24.175 9.545 ;
        RECT 23.195 9.360 24.175 9.500 ;
        RECT 23.195 9.315 23.485 9.360 ;
        RECT 23.885 9.315 24.175 9.360 ;
      LAYER met2 ;
        RECT 23.550 11.680 23.830 13.680 ;
        RECT 23.620 10.015 23.760 11.680 ;
        RECT 23.900 10.015 24.220 10.075 ;
        RECT 23.620 9.875 24.220 10.015 ;
        RECT 23.900 9.815 24.220 9.875 ;
    END
  END gpio_defaults[29]
  PIN gpio_defaults[30]
    PORT
      LAYER li1 ;
        RECT 25.155 3.635 25.675 5.185 ;
      LAYER met1 ;
        RECT 24.575 3.980 24.865 4.025 ;
        RECT 25.265 3.980 25.555 4.025 ;
        RECT 24.575 3.840 25.555 3.980 ;
        RECT 24.575 3.795 24.865 3.840 ;
        RECT 25.265 3.795 25.555 3.840 ;
        RECT 25.355 3.555 25.495 3.795 ;
        RECT 25.310 3.235 25.570 3.555 ;
      LAYER met2 ;
        RECT 25.280 3.465 25.600 3.525 ;
        RECT 25.000 3.325 25.600 3.465 ;
        RECT 25.000 2.000 25.140 3.325 ;
        RECT 25.280 3.265 25.600 3.325 ;
        RECT 24.930 0.000 25.210 2.000 ;
    END
  END gpio_defaults[30]
  PIN gpio_defaults[31]
    PORT
      LAYER li1 ;
        RECT 25.155 9.075 25.675 10.625 ;
      LAYER met1 ;
        RECT 25.310 9.785 25.570 10.105 ;
        RECT 25.355 9.545 25.495 9.785 ;
        RECT 24.575 9.500 24.865 9.545 ;
        RECT 25.265 9.500 25.555 9.545 ;
        RECT 24.575 9.360 25.555 9.500 ;
        RECT 24.575 9.315 24.865 9.360 ;
        RECT 25.265 9.315 25.555 9.360 ;
      LAYER met2 ;
        RECT 24.930 11.680 25.210 13.680 ;
        RECT 25.000 10.015 25.140 11.680 ;
        RECT 25.280 10.015 25.600 10.075 ;
        RECT 25.000 9.875 25.600 10.015 ;
        RECT 25.280 9.815 25.600 9.875 ;
    END
  END gpio_defaults[31]
  OBS
      LAYER pwell ;
        RECT 0.005 8.265 1.375 9.075 ;
        RECT 25.765 8.265 27.135 9.075 ;
        RECT 0.145 8.055 0.315 8.265 ;
        RECT 1.525 8.215 1.695 8.245 ;
        RECT 1.520 8.105 1.695 8.215 ;
        RECT 1.525 8.055 1.695 8.105 ;
        RECT 1.985 8.075 2.155 8.245 ;
        RECT 3.365 8.075 3.535 8.245 ;
        RECT 4.285 8.055 4.455 8.245 ;
        RECT 4.745 8.075 4.915 8.245 ;
        RECT 6.125 8.075 6.295 8.245 ;
        RECT 7.505 8.075 7.675 8.245 ;
        RECT 8.885 8.075 9.055 8.245 ;
        RECT 9.805 8.055 9.975 8.245 ;
        RECT 10.720 8.105 10.840 8.215 ;
        RECT 11.185 8.075 11.355 8.245 ;
        RECT 12.565 8.075 12.735 8.245 ;
        RECT 13.945 8.075 14.115 8.245 ;
        RECT 15.325 8.215 15.495 8.245 ;
        RECT 15.320 8.105 15.495 8.215 ;
        RECT 15.325 8.055 15.495 8.105 ;
        RECT 15.785 8.075 15.955 8.245 ;
        RECT 17.165 8.075 17.335 8.245 ;
        RECT 18.545 8.075 18.715 8.245 ;
        RECT 19.925 8.075 20.095 8.245 ;
        RECT 20.845 8.055 21.015 8.245 ;
        RECT 21.305 8.075 21.475 8.245 ;
        RECT 22.680 8.105 22.800 8.215 ;
        RECT 23.145 8.075 23.315 8.245 ;
        RECT 23.605 8.055 23.775 8.245 ;
        RECT 24.525 8.075 24.695 8.245 ;
        RECT 25.440 8.105 25.560 8.215 ;
        RECT 26.825 8.055 26.995 8.265 ;
        RECT 0.005 7.245 1.375 8.055 ;
        RECT 1.385 7.245 4.135 8.055 ;
        RECT 4.145 7.245 9.655 8.055 ;
        RECT 9.665 7.245 15.175 8.055 ;
        RECT 15.185 7.245 20.695 8.055 ;
        RECT 20.705 7.245 22.535 8.055 ;
        RECT 23.465 7.245 25.295 8.055 ;
        RECT 25.765 7.245 27.135 8.055 ;
        RECT 0.005 2.825 1.375 3.635 ;
        RECT 25.765 2.825 27.135 3.635 ;
        RECT 0.145 2.635 0.315 2.825 ;
        RECT 1.520 2.665 1.640 2.775 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 10.720 2.665 10.840 2.775 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 15.320 2.665 15.440 2.775 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 17.165 2.635 17.335 2.805 ;
        RECT 18.545 2.635 18.715 2.805 ;
        RECT 19.925 2.635 20.095 2.805 ;
        RECT 21.305 2.635 21.475 2.805 ;
        RECT 23.145 2.635 23.315 2.805 ;
        RECT 24.525 2.635 24.695 2.805 ;
        RECT 26.825 2.635 26.995 2.825 ;
      LAYER li1 ;
        RECT 1.925 8.415 2.445 9.900 ;
        RECT 3.305 8.415 3.825 9.900 ;
        RECT 4.685 8.415 5.205 9.900 ;
        RECT 6.065 8.415 6.585 9.900 ;
        RECT 7.445 8.415 7.965 9.900 ;
        RECT 8.825 8.415 9.345 9.900 ;
        RECT 11.125 8.415 11.645 9.900 ;
        RECT 12.505 8.415 13.025 9.900 ;
        RECT 13.885 8.415 14.405 9.900 ;
        RECT 15.725 8.415 16.245 9.900 ;
        RECT 17.105 8.415 17.625 9.900 ;
        RECT 18.485 8.415 19.005 9.900 ;
        RECT 19.865 8.415 20.385 9.900 ;
        RECT 21.245 8.415 21.765 9.900 ;
        RECT 23.085 8.415 23.605 9.900 ;
        RECT 24.465 8.415 24.985 9.900 ;
        RECT 1.925 2.975 2.445 4.460 ;
        RECT 3.305 2.975 3.825 4.460 ;
        RECT 4.685 2.975 5.205 4.460 ;
        RECT 6.065 2.975 6.585 4.460 ;
        RECT 7.445 2.975 7.965 4.460 ;
        RECT 8.825 2.975 9.345 4.460 ;
        RECT 11.125 2.975 11.645 4.460 ;
        RECT 12.505 2.975 13.025 4.460 ;
        RECT 13.885 2.975 14.405 4.460 ;
        RECT 15.725 2.975 16.245 4.460 ;
        RECT 17.105 2.975 17.625 4.460 ;
        RECT 18.485 2.975 19.005 4.460 ;
        RECT 19.865 2.975 20.385 4.460 ;
        RECT 21.245 2.975 21.765 4.460 ;
        RECT 23.085 2.975 23.605 4.460 ;
        RECT 24.465 2.975 24.985 4.460 ;
  END
END project_id_rom_32bit
END LIBRARY

