VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_QSPI_XIP_CTRL_AHBL
  CLASS BLOCK ;
  FOREIGN EF_QSPI_XIP_CTRL_AHBL ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 500.000 ;
  PIN HADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 496.000 41.310 500.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 151.430 496.000 151.710 500.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.470 496.000 162.750 500.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.510 496.000 173.790 500.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 184.550 496.000 184.830 500.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.590 496.000 195.870 500.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.630 496.000 206.910 500.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.670 496.000 217.950 500.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 228.710 496.000 228.990 500.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 239.750 496.000 240.030 500.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 250.790 496.000 251.070 500.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 496.000 52.350 500.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 261.830 496.000 262.110 500.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 272.870 496.000 273.150 500.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.910 496.000 284.190 500.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 294.950 496.000 295.230 500.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 496.000 306.270 500.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 496.000 317.310 500.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 496.000 328.350 500.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 496.000 339.390 500.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 496.000 350.430 500.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 496.000 361.470 500.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 63.110 496.000 63.390 500.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 496.000 372.510 500.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 496.000 383.550 500.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.150 496.000 74.430 500.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 85.190 496.000 85.470 500.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.563400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 96.230 496.000 96.510 500.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.276700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 107.270 496.000 107.550 500.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.177200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 118.310 496.000 118.590 500.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.276700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 129.350 496.000 129.630 500.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 140.390 496.000 140.670 500.000 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 7.910 496.000 8.190 500.000 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 449.510 496.000 449.790 500.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 559.910 496.000 560.190 500.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 570.950 496.000 571.230 500.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 581.990 496.000 582.270 500.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 593.030 496.000 593.310 500.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 604.070 496.000 604.350 500.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 615.110 496.000 615.390 500.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 626.150 496.000 626.430 500.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 637.190 496.000 637.470 500.000 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 648.230 496.000 648.510 500.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 659.270 496.000 659.550 500.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 460.550 496.000 460.830 500.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 670.310 496.000 670.590 500.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 681.350 496.000 681.630 500.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 692.390 496.000 692.670 500.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 703.430 496.000 703.710 500.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 714.470 496.000 714.750 500.000 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 725.510 496.000 725.790 500.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 736.550 496.000 736.830 500.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 747.590 496.000 747.870 500.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 758.630 496.000 758.910 500.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 769.670 496.000 769.950 500.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 471.590 496.000 471.870 500.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 780.710 496.000 780.990 500.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 791.750 496.000 792.030 500.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 482.630 496.000 482.910 500.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 493.670 496.000 493.950 500.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 504.710 496.000 504.990 500.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 515.750 496.000 516.030 500.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 526.790 496.000 527.070 500.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 537.830 496.000 538.110 500.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 548.870 496.000 549.150 500.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 427.430 496.000 427.710 500.000 ;
    END
  END HREADY
  PIN HREADYOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 438.470 496.000 438.750 500.000 ;
    END
  END HREADYOUT
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 18.950 496.000 19.230 500.000 ;
    END
  END HRESETn
  PIN HSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.990 496.000 30.270 500.000 ;
    END
  END HSEL
  PIN HTRANS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 496.000 394.590 500.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 405.350 496.000 405.630 500.000 ;
    END
  END HTRANS[1]
  PIN HWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 496.000 416.670 500.000 ;
    END
  END HWRITE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.340 10.640 105.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.340 10.640 185.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.340 10.640 265.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.340 10.640 345.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 10.640 425.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.340 10.640 505.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 584.340 10.640 585.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.340 10.640 665.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.340 10.640 745.940 487.120 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.040 10.640 102.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.040 10.640 182.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.040 10.640 342.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 581.040 10.640 582.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.040 10.640 662.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 487.120 ;
    END
  END VPWR
  PIN ce_n
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END ce_n
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END din[0]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END din[1]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END din[2]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END din[3]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END dout[1]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END dout[2]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END dout[3]
  PIN douten[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END douten[0]
  PIN douten[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END douten[1]
  PIN douten[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END douten[2]
  PIN douten[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END douten[3]
  PIN sck
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END sck
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 794.610 487.070 ;
      LAYER li1 ;
        RECT 5.520 10.795 794.420 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 794.420 497.040 ;
      LAYER met2 ;
        RECT 8.470 495.720 18.670 497.070 ;
        RECT 19.510 495.720 29.710 497.070 ;
        RECT 30.550 495.720 40.750 497.070 ;
        RECT 41.590 495.720 51.790 497.070 ;
        RECT 52.630 495.720 62.830 497.070 ;
        RECT 63.670 495.720 73.870 497.070 ;
        RECT 74.710 495.720 84.910 497.070 ;
        RECT 85.750 495.720 95.950 497.070 ;
        RECT 96.790 495.720 106.990 497.070 ;
        RECT 107.830 495.720 118.030 497.070 ;
        RECT 118.870 495.720 129.070 497.070 ;
        RECT 129.910 495.720 140.110 497.070 ;
        RECT 140.950 495.720 151.150 497.070 ;
        RECT 151.990 495.720 162.190 497.070 ;
        RECT 163.030 495.720 173.230 497.070 ;
        RECT 174.070 495.720 184.270 497.070 ;
        RECT 185.110 495.720 195.310 497.070 ;
        RECT 196.150 495.720 206.350 497.070 ;
        RECT 207.190 495.720 217.390 497.070 ;
        RECT 218.230 495.720 228.430 497.070 ;
        RECT 229.270 495.720 239.470 497.070 ;
        RECT 240.310 495.720 250.510 497.070 ;
        RECT 251.350 495.720 261.550 497.070 ;
        RECT 262.390 495.720 272.590 497.070 ;
        RECT 273.430 495.720 283.630 497.070 ;
        RECT 284.470 495.720 294.670 497.070 ;
        RECT 295.510 495.720 305.710 497.070 ;
        RECT 306.550 495.720 316.750 497.070 ;
        RECT 317.590 495.720 327.790 497.070 ;
        RECT 328.630 495.720 338.830 497.070 ;
        RECT 339.670 495.720 349.870 497.070 ;
        RECT 350.710 495.720 360.910 497.070 ;
        RECT 361.750 495.720 371.950 497.070 ;
        RECT 372.790 495.720 382.990 497.070 ;
        RECT 383.830 495.720 394.030 497.070 ;
        RECT 394.870 495.720 405.070 497.070 ;
        RECT 405.910 495.720 416.110 497.070 ;
        RECT 416.950 495.720 427.150 497.070 ;
        RECT 427.990 495.720 438.190 497.070 ;
        RECT 439.030 495.720 449.230 497.070 ;
        RECT 450.070 495.720 460.270 497.070 ;
        RECT 461.110 495.720 471.310 497.070 ;
        RECT 472.150 495.720 482.350 497.070 ;
        RECT 483.190 495.720 493.390 497.070 ;
        RECT 494.230 495.720 504.430 497.070 ;
        RECT 505.270 495.720 515.470 497.070 ;
        RECT 516.310 495.720 526.510 497.070 ;
        RECT 527.350 495.720 537.550 497.070 ;
        RECT 538.390 495.720 548.590 497.070 ;
        RECT 549.430 495.720 559.630 497.070 ;
        RECT 560.470 495.720 570.670 497.070 ;
        RECT 571.510 495.720 581.710 497.070 ;
        RECT 582.550 495.720 592.750 497.070 ;
        RECT 593.590 495.720 603.790 497.070 ;
        RECT 604.630 495.720 614.830 497.070 ;
        RECT 615.670 495.720 625.870 497.070 ;
        RECT 626.710 495.720 636.910 497.070 ;
        RECT 637.750 495.720 647.950 497.070 ;
        RECT 648.790 495.720 658.990 497.070 ;
        RECT 659.830 495.720 670.030 497.070 ;
        RECT 670.870 495.720 681.070 497.070 ;
        RECT 681.910 495.720 692.110 497.070 ;
        RECT 692.950 495.720 703.150 497.070 ;
        RECT 703.990 495.720 714.190 497.070 ;
        RECT 715.030 495.720 725.230 497.070 ;
        RECT 726.070 495.720 736.270 497.070 ;
        RECT 737.110 495.720 747.310 497.070 ;
        RECT 748.150 495.720 758.350 497.070 ;
        RECT 759.190 495.720 769.390 497.070 ;
        RECT 770.230 495.720 780.430 497.070 ;
        RECT 781.270 495.720 791.470 497.070 ;
        RECT 792.310 495.720 792.940 497.070 ;
        RECT 7.920 4.280 792.940 495.720 ;
        RECT 7.920 4.000 28.790 4.280 ;
        RECT 29.630 4.000 85.830 4.280 ;
        RECT 86.670 4.000 142.870 4.280 ;
        RECT 143.710 4.000 199.910 4.280 ;
        RECT 200.750 4.000 256.950 4.280 ;
        RECT 257.790 4.000 313.990 4.280 ;
        RECT 314.830 4.000 371.030 4.280 ;
        RECT 371.870 4.000 428.070 4.280 ;
        RECT 428.910 4.000 485.110 4.280 ;
        RECT 485.950 4.000 542.150 4.280 ;
        RECT 542.990 4.000 599.190 4.280 ;
        RECT 600.030 4.000 656.230 4.280 ;
        RECT 657.070 4.000 713.270 4.280 ;
        RECT 714.110 4.000 770.310 4.280 ;
        RECT 771.150 4.000 792.940 4.280 ;
      LAYER met3 ;
        RECT 16.165 10.715 789.755 487.045 ;
      LAYER met4 ;
        RECT 23.295 18.535 23.940 486.025 ;
        RECT 26.340 18.535 100.640 486.025 ;
        RECT 103.040 18.535 103.940 486.025 ;
        RECT 106.340 18.535 180.640 486.025 ;
        RECT 183.040 18.535 183.940 486.025 ;
        RECT 186.340 18.535 260.640 486.025 ;
        RECT 263.040 18.535 263.940 486.025 ;
        RECT 266.340 18.535 340.640 486.025 ;
        RECT 343.040 18.535 343.940 486.025 ;
        RECT 346.340 18.535 420.640 486.025 ;
        RECT 423.040 18.535 423.940 486.025 ;
        RECT 426.340 18.535 500.640 486.025 ;
        RECT 503.040 18.535 503.940 486.025 ;
        RECT 506.340 18.535 580.640 486.025 ;
        RECT 583.040 18.535 583.940 486.025 ;
        RECT 586.340 18.535 660.640 486.025 ;
        RECT 663.040 18.535 663.940 486.025 ;
        RECT 666.340 18.535 740.640 486.025 ;
        RECT 743.040 18.535 743.940 486.025 ;
        RECT 746.340 18.535 749.505 486.025 ;
  END
END EF_QSPI_XIP_CTRL_AHBL
END LIBRARY

