magic
tech sky130A
magscale 1 2
timestamp 1581648494
<< checkpaint >>
rect -1251 -1260 719153 1039064
use frigate_core  frigate_core_0
timestamp 1581648494
transform 1 0 41151 0 1 41204
box -700 -698 636300 956576
use panamax  panamax_0
timestamp 1581648494
transform 1 0 151 0 1 204
box -142 -204 717742 1037600
<< labels >>
flabel metal5 s 704908 870904 704908 870904 0 FreeSans 37500 0 0 0 gpio2_4
flabel metal5 s 704908 891904 704908 891904 0 FreeSans 37500 0 0 0 gpio2_5
flabel metal5 s 704908 912904 704908 912904 0 FreeSans 37500 0 0 0 gpio2_6
flabel metal5 s 704908 933904 704908 933904 0 FreeSans 37500 0 0 0 gpio2_7
flabel metal5 s 704831 954904 704831 954904 0 FreeSans 37500 0 0 0 vccd1_1
flabel metal5 s 704831 978904 704831 978904 0 FreeSans 37500 0 0 0 vddio_3
flabel metal5 s 704831 530904 704831 530904 0 FreeSans 37500 0 0 0 vssio_1
flabel metal5 s 705247 560538 705247 560538 0 FreeSans 37500 0 0 0 gpio1_4
flabel metal5 s 705247 593538 705247 593538 0 FreeSans 37500 0 0 0 gpio1_5
flabel metal5 s 705247 626538 705247 626538 0 FreeSans 37500 0 0 0 gpio1_6
flabel metal5 s 705247 659538 705247 659538 0 FreeSans 37500 0 0 0 gpio1_7
flabel metal5 s 704908 870904 704908 870904 0 FreeSans 37500 0 0 0 gpio2_4
flabel metal5 s 704908 891904 704908 891904 0 FreeSans 37500 0 0 0 gpio2_5
flabel metal5 s 704908 912904 704908 912904 0 FreeSans 37500 0 0 0 gpio2_6
flabel metal5 s 704908 933904 704908 933904 0 FreeSans 37500 0 0 0 gpio2_7
flabel metal5 s 704831 954904 704831 954904 0 FreeSans 37500 0 0 0 vccd1_1
flabel metal5 s 704831 682904 704831 682904 0 FreeSans 37500 0 0 0 vddio_2
flabel metal5 s 704831 702904 704831 702904 0 FreeSans 37500 0 0 0 vdda1_1
flabel metal5 s 704831 726904 704831 726904 0 FreeSans 37500 0 0 0 vssa1_1
flabel metal5 s 704831 746904 704831 746904 0 FreeSans 37500 0 0 0 vssd1_1
flabel metal5 s 704908 766904 704908 766904 0 FreeSans 37500 0 0 0 gpio2_0
flabel metal5 s 704908 787904 704908 787904 0 FreeSans 37500 0 0 0 gpio2_1
flabel metal5 s 704908 808904 704908 808904 0 FreeSans 37500 0 0 0 gpio2_2
flabel metal5 s 704908 829904 704908 829904 0 FreeSans 37500 0 0 0 gpio2_3
flabel metal5 s 704831 850904 704831 850904 0 FreeSans 37500 0 0 0 vssio_2
flabel metal5 s 704908 870904 704908 870904 0 FreeSans 37500 0 0 0 gpio2_4
flabel metal5 s 704908 891904 704908 891904 0 FreeSans 37500 0 0 0 gpio2_5
flabel metal5 s 704908 912904 704908 912904 0 FreeSans 37500 0 0 0 gpio2_6
flabel metal5 s 704908 933904 704908 933904 0 FreeSans 37500 0 0 0 gpio2_7
flabel metal5 s 704831 954904 704831 954904 0 FreeSans 37500 0 0 0 vccd1_1
flabel metal5 s 359451 1024884 359451 1024884 0 FreeSans 37500 0 0 0 analog_0
flabel metal5 s 382451 1024884 382451 1024884 0 FreeSans 37500 0 0 0 vdda0_0
flabel metal5 s 405451 1024884 405451 1024884 0 FreeSans 37500 0 0 0 vddio_4
flabel metal5 s 429451 1024961 429451 1024961 0 FreeSans 37500 0 0 0 gpio3_7
flabel metal5 s 453451 1024961 453451 1024961 0 FreeSans 37500 0 0 0 gpio3_6
flabel metal5 s 477451 1024961 477451 1024961 0 FreeSans 37500 0 0 0 gpio3_5
flabel metal5 s 501451 1024961 501451 1024961 0 FreeSans 37500 0 0 0 gpio3_4
flabel metal5 s 524451 1024884 524451 1024884 0 FreeSans 37500 0 0 0 vccd1_2
flabel metal5 s 547451 1024884 547451 1024884 0 FreeSans 37500 0 0 0 vssio_3
flabel metal5 s 571451 1024961 571451 1024961 0 FreeSans 37500 0 0 0 gpio3_3
flabel metal5 s 595451 1024961 595451 1024961 0 FreeSans 37500 0 0 0 gpio3_2
flabel metal5 s 619451 1024961 619451 1024961 0 FreeSans 37500 0 0 0 gpio3_1
flabel metal5 s 643451 1024961 643451 1024961 0 FreeSans 37500 0 0 0 gpio3_0
flabel metal5 s 666451 1024884 666451 1024884 0 FreeSans 37500 0 0 0 vssd1_2
flabel metal5 s 76451 1024961 76451 1024961 0 FreeSans 37500 0 0 0 gpio4_7
flabel metal5 s 100451 1024961 100451 1024961 0 FreeSans 37500 0 0 0 gpio4_6
flabel metal5 s 124451 1024961 124451 1024961 0 FreeSans 37500 0 0 0 gpio4_5
flabel metal5 s 148451 1024961 148451 1024961 0 FreeSans 37500 0 0 0 gpio4_4
flabel metal5 s 171451 1024884 171451 1024884 0 FreeSans 37500 0 0 0 vssio_4
flabel metal5 s 194451 1024884 194451 1024884 0 FreeSans 37500 0 0 0 vssd2_0
flabel metal5 s 218451 1024961 218451 1024961 0 FreeSans 37500 0 0 0 gpio4_3
flabel metal5 s 242451 1024961 242451 1024961 0 FreeSans 37500 0 0 0 gpio4_2
flabel metal5 s 266451 1024961 266451 1024961 0 FreeSans 37500 0 0 0 gpio4_1
flabel metal5 s 290451 1024961 290451 1024961 0 FreeSans 37500 0 0 0 gpio4_0
flabel metal5 s 313451 1024884 313451 1024884 0 FreeSans 37500 0 0 0 vssa0_0
flabel metal5 s 336451 1024884 336451 1024884 0 FreeSans 37500 0 0 0 analog_1
flabel metal5 s 52451 1024884 52451 1024884 0 FreeSans 37500 0 0 0 vccd2_0
flabel metal5 s 13071 533704 13071 533704 0 FreeSans 37500 0 0 0 vssio_6
flabel metal5 s 12655 557070 12655 557070 0 FreeSans 37500 0 0 0 gpio6_3
flabel metal5 s 12655 590070 12655 590070 0 FreeSans 37500 0 0 0 gpio6_2
flabel metal5 s 12655 623070 12655 623070 0 FreeSans 37500 0 0 0 gpio6_1
flabel metal5 s 12655 656070 12655 656070 0 FreeSans 37500 0 0 0 gpio6_0
flabel metal5 s 13071 685704 13071 685704 0 FreeSans 37500 0 0 0 vddio_6
flabel metal5 s 13071 705704 13071 705704 0 FreeSans 37500 0 0 0 vdda2_0
flabel metal5 s 13071 728704 13071 728704 0 FreeSans 37500 0 0 0 vssa2_0
flabel metal5 s 13071 748704 13071 748704 0 FreeSans 37500 0 0 0 vccd2_1
flabel metal5 s 12994 769704 12994 769704 0 FreeSans 37500 0 0 0 gpio5_7
flabel metal5 s 12994 790704 12994 790704 0 FreeSans 37500 0 0 0 gpio5_6
flabel metal5 s 12994 811704 12994 811704 0 FreeSans 37500 0 0 0 gpio5_5
flabel metal5 s 12994 832704 12994 832704 0 FreeSans 37500 0 0 0 gpio5_4
flabel metal5 s 13071 852704 13071 852704 0 FreeSans 37500 0 0 0 vssio_5
flabel metal5 s 12994 873704 12994 873704 0 FreeSans 37500 0 0 0 gpio5_3
flabel metal5 s 12994 894704 12994 894704 0 FreeSans 37500 0 0 0 gpio5_2
flabel metal5 s 12994 915704 12994 915704 0 FreeSans 37500 0 0 0 gpio5_1
flabel metal5 s 12994 936704 12994 936704 0 FreeSans 37500 0 0 0 gpio5_0
flabel metal5 s 13071 956704 13071 956704 0 FreeSans 37500 0 0 0 vssd2_1
flabel metal5 s 13071 979704 13071 979704 0 FreeSans 37500 0 0 0 vddio_5
flabel metal5 s 13071 190104 13071 190104 0 FreeSans 37500 0 0 0 vssio_7
flabel metal5 s 12994 211104 12994 211104 0 FreeSans 37500 0 0 0 gpio7_3
flabel metal5 s 12994 232104 12994 232104 0 FreeSans 37500 0 0 0 gpio7_2
flabel metal5 s 12994 253104 12994 253104 0 FreeSans 37500 0 0 0 gpio7_1
flabel metal5 s 12994 274104 12994 274104 0 FreeSans 37500 0 0 0 gpio7_0
flabel metal5 s 13071 294104 13071 294104 0 FreeSans 37500 0 0 0 vddio_7
flabel metal5 s 13071 314104 13071 314104 0 FreeSans 37500 0 0 0 vdda2_1
flabel metal5 s 13071 337104 13071 337104 0 FreeSans 37500 0 0 0 vssa2_1
flabel metal5 s 12655 360470 12655 360470 0 FreeSans 37500 0 0 0 gpio6_7
flabel metal5 s 12655 393470 12655 393470 0 FreeSans 37500 0 0 0 gpio6_6
flabel metal5 s 12655 426470 12655 426470 0 FreeSans 37500 0 0 0 gpio6_5
flabel metal5 s 12655 459470 12655 459470 0 FreeSans 37500 0 0 0 gpio6_4
flabel metal5 s 13071 489104 13071 489104 0 FreeSans 37500 0 0 0 vssd2_2
flabel metal5 s 13071 63104 13071 63104 0 FreeSans 37500 0 0 0 vddio_8
flabel metal5 s 12994 84104 12994 84104 0 FreeSans 37500 0 0 0 gpio7_7
flabel metal5 s 12994 105104 12994 105104 0 FreeSans 37500 0 0 0 gpio7_6
flabel metal5 s 12994 126104 12994 126104 0 FreeSans 37500 0 0 0 gpio7_5
flabel metal5 s 12994 147104 12994 147104 0 FreeSans 37500 0 0 0 gpio7_4
flabel metal5 s 13071 167104 13071 167104 0 FreeSans 37500 0 0 0 vccd2_2
flabel metal5 s 167651 13047 167651 13047 0 FreeSans 37500 0 0 0 gpio8_2
flabel metal5 s 190651 13047 190651 13047 0 FreeSans 37500 0 0 0 gpio8_3
flabel metal5 s 213651 13124 213651 13124 0 FreeSans 37500 0 0 0 vssio_8
flabel metal5 s 235651 13124 235651 13124 0 FreeSans 37500 0 0 0 vssd0_0
flabel metal5 s 257651 13124 257651 13124 0 FreeSans 37500 0 0 0 xi0
flabel metal5 s 279651 13124 279651 13124 0 FreeSans 37500 0 0 0 xo0
flabel metal5 s 301651 13124 301651 13124 0 FreeSans 37500 0 0 0 xi1
flabel metal5 s 323651 13124 323651 13124 0 FreeSans 37500 0 0 0 xo1
flabel metal5 s 345651 13124 345651 13124 0 FreeSans 37500 0 0 0 vddio_9
flabel metal5 s 54651 13124 54651 13124 0 FreeSans 37500 0 0 0 vccd0_0
flabel metal5 s 76651 13047 76651 13047 0 FreeSans 37500 0 0 0 select
flabel metal5 s 99651 13124 99651 13124 0 FreeSans 37500 0 0 0 resetb
flabel metal5 s 121651 13047 121651 13047 0 FreeSans 37500 0 0 0 gpio8_0
flabel metal5 s 144651 13047 144651 13047 0 FreeSans 37500 0 0 0 gpio8_1
flabel metal5 s 704908 248304 704908 248304 0 FreeSans 37500 0 0 0 gpio0_6
flabel metal5 s 704908 269304 704908 269304 0 FreeSans 37500 0 0 0 gpio0_7
flabel metal5 s 704831 290304 704831 290304 0 FreeSans 37500 0 0 0 vddio_1
flabel metal5 s 704831 334304 704831 334304 0 FreeSans 37500 0 0 0 vssa1_0
flabel metal5 s 705247 363938 705247 363938 0 FreeSans 37500 0 0 0 gpio1_0
flabel metal5 s 704831 310304 704831 310304 0 FreeSans 37500 0 0 0 vdda1_0
flabel metal5 s 705247 396938 705247 396938 0 FreeSans 37500 0 0 0 gpio1_1
flabel metal5 s 705247 429938 705247 429938 0 FreeSans 37500 0 0 0 gpio1_2
flabel metal5 s 705247 462938 705247 462938 0 FreeSans 37500 0 0 0 gpio1_3
flabel metal5 s 704831 486304 704831 486304 0 FreeSans 37500 0 0 0 vccd1_0
flabel metal5 s 704831 186304 704831 186304 0 FreeSans 37500 0 0 0 vssio_0
flabel metal5 s 704908 206304 704908 206304 0 FreeSans 37500 0 0 0 gpio0_4
flabel metal5 s 704908 227304 704908 227304 0 FreeSans 37500 0 0 0 gpio0_5
flabel metal5 s 704831 62304 704831 62304 0 FreeSans 37500 0 0 0 vddio_0
flabel metal5 s 704908 82304 704908 82304 0 FreeSans 37500 0 0 0 gpio0_0
flabel metal5 s 704908 103304 704908 103304 0 FreeSans 37500 0 0 0 gpio0_1
flabel metal5 s 704908 124304 704908 124304 0 FreeSans 37500 0 0 0 gpio0_2
flabel metal5 s 704908 145304 704908 145304 0 FreeSans 37500 0 0 0 gpio0_3
flabel metal5 s 704831 166304 704831 166304 0 FreeSans 37500 0 0 0 vssd1_0
flabel metal5 s 371651 13124 371651 13124 0 FreeSans 37500 0 0 0 vccd0_1
flabel metal5 s 393651 13047 393651 13047 0 FreeSans 37500 0 0 0 gpio8_4
flabel metal5 s 416651 13047 416651 13047 0 FreeSans 37500 0 0 0 gpio8_5
flabel metal5 s 439651 13047 439651 13047 0 FreeSans 37500 0 0 0 gpio8_6
flabel metal5 s 462651 13047 462651 13047 0 FreeSans 37500 0 0 0 gpio8_7
flabel metal5 s 485651 13124 485651 13124 0 FreeSans 37500 0 0 0 vssio_9
flabel metal5 s 507651 13124 507651 13124 0 FreeSans 37500 0 0 0 vssa3_0
flabel metal5 s 533651 13124 533651 13124 0 FreeSans 37500 0 0 0 vdda3_0
flabel metal5 s 559651 13124 559651 13124 0 FreeSans 37500 0 0 0 vssd0_1
flabel metal5 s 619848 18272 619848 18272 0 FreeSans 37500 0 0 0 sio0
flabel metal5 s 642453 18272 642453 18272 0 FreeSans 37500 0 0 0 sio1
<< end >>
