VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ctu_can
  CLASS BLOCK ;
  FOREIGN ctu_can ;
  ORIGIN 0.000 0.000 ;
  SIZE 580.000 BY 580.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.340 10.640 105.940 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.340 10.640 185.940 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.340 10.640 265.940 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.340 10.640 345.940 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 10.640 425.940 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.340 10.640 505.940 568.720 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.040 10.640 102.640 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.040 10.640 182.640 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.040 10.640 342.640 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 568.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 568.720 ;
    END
  END VPWR
  PIN adress[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 576.000 457.000 580.000 457.600 ;
    END
  END adress[0]
  PIN adress[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 484.200 580.000 484.800 ;
    END
  END adress[10]
  PIN adress[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 486.920 580.000 487.520 ;
    END
  END adress[11]
  PIN adress[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 576.000 489.640 580.000 490.240 ;
    END
  END adress[12]
  PIN adress[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 576.000 492.360 580.000 492.960 ;
    END
  END adress[13]
  PIN adress[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 576.000 495.080 580.000 495.680 ;
    END
  END adress[14]
  PIN adress[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 576.000 497.800 580.000 498.400 ;
    END
  END adress[15]
  PIN adress[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 576.000 459.720 580.000 460.320 ;
    END
  END adress[1]
  PIN adress[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 462.440 580.000 463.040 ;
    END
  END adress[2]
  PIN adress[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 465.160 580.000 465.760 ;
    END
  END adress[3]
  PIN adress[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 467.880 580.000 468.480 ;
    END
  END adress[4]
  PIN adress[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 470.600 580.000 471.200 ;
    END
  END adress[5]
  PIN adress[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 473.320 580.000 473.920 ;
    END
  END adress[6]
  PIN adress[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 476.040 580.000 476.640 ;
    END
  END adress[7]
  PIN adress[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 478.760 580.000 479.360 ;
    END
  END adress[8]
  PIN adress[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 481.480 580.000 482.080 ;
    END
  END adress[9]
  PIN can_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 14.810 576.000 15.090 580.000 ;
    END
  END can_rx
  PIN can_tx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 35.970 576.000 36.250 580.000 ;
    END
  END can_tx
  PIN clk_sys
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 84.360 580.000 84.960 ;
    END
  END clk_sys
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 89.800 580.000 90.400 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 117.000 580.000 117.600 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 119.720 580.000 120.320 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 122.440 580.000 123.040 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 125.160 580.000 125.760 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 127.880 580.000 128.480 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 130.600 580.000 131.200 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 133.320 580.000 133.920 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 136.040 580.000 136.640 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 138.760 580.000 139.360 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 141.480 580.000 142.080 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 92.520 580.000 93.120 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 144.200 580.000 144.800 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 146.920 580.000 147.520 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 149.640 580.000 150.240 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 152.360 580.000 152.960 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 155.080 580.000 155.680 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 157.800 580.000 158.400 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 160.520 580.000 161.120 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 163.240 580.000 163.840 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 165.960 580.000 166.560 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 168.680 580.000 169.280 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 95.240 580.000 95.840 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 171.400 580.000 172.000 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 174.120 580.000 174.720 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 97.960 580.000 98.560 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 100.680 580.000 101.280 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 103.400 580.000 104.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 106.120 580.000 106.720 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 108.840 580.000 109.440 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 111.560 580.000 112.160 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 114.280 580.000 114.880 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 369.960 580.000 370.560 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 397.160 580.000 397.760 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 399.880 580.000 400.480 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 402.600 580.000 403.200 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 405.320 580.000 405.920 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 408.040 580.000 408.640 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 410.760 580.000 411.360 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 413.480 580.000 414.080 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 416.200 580.000 416.800 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 418.920 580.000 419.520 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 421.640 580.000 422.240 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 372.680 580.000 373.280 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 424.360 580.000 424.960 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 427.080 580.000 427.680 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 429.800 580.000 430.400 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 432.520 580.000 433.120 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 435.240 580.000 435.840 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 437.960 580.000 438.560 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 440.680 580.000 441.280 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 443.400 580.000 444.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 446.120 580.000 446.720 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 448.840 580.000 449.440 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 375.400 580.000 376.000 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 451.560 580.000 452.160 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 454.280 580.000 454.880 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 378.120 580.000 378.720 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 380.840 580.000 381.440 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 383.560 580.000 384.160 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 386.280 580.000 386.880 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 389.000 580.000 389.600 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 391.720 580.000 392.320 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 394.440 580.000 395.040 ;
    END
  END data_out[9]
  PIN int_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 81.640 580.000 82.240 ;
    END
  END int_
  PIN res_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 87.080 580.000 87.680 ;
    END
  END res_n
  PIN sbe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 176.840 580.000 177.440 ;
    END
  END sbe[0]
  PIN sbe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 179.560 580.000 180.160 ;
    END
  END sbe[1]
  PIN sbe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 182.280 580.000 182.880 ;
    END
  END sbe[2]
  PIN sbe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 185.000 580.000 185.600 ;
    END
  END sbe[3]
  PIN scs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 187.720 580.000 188.320 ;
    END
  END scs
  PIN srd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 190.440 580.000 191.040 ;
    END
  END srd
  PIN swr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 193.160 580.000 193.760 ;
    END
  END swr
  PIN timestamp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 195.880 580.000 196.480 ;
    END
  END timestamp[0]
  PIN timestamp[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 223.080 580.000 223.680 ;
    END
  END timestamp[10]
  PIN timestamp[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 225.800 580.000 226.400 ;
    END
  END timestamp[11]
  PIN timestamp[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 228.520 580.000 229.120 ;
    END
  END timestamp[12]
  PIN timestamp[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 231.240 580.000 231.840 ;
    END
  END timestamp[13]
  PIN timestamp[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 233.960 580.000 234.560 ;
    END
  END timestamp[14]
  PIN timestamp[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 236.680 580.000 237.280 ;
    END
  END timestamp[15]
  PIN timestamp[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 239.400 580.000 240.000 ;
    END
  END timestamp[16]
  PIN timestamp[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 242.120 580.000 242.720 ;
    END
  END timestamp[17]
  PIN timestamp[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 244.840 580.000 245.440 ;
    END
  END timestamp[18]
  PIN timestamp[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 247.560 580.000 248.160 ;
    END
  END timestamp[19]
  PIN timestamp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 198.600 580.000 199.200 ;
    END
  END timestamp[1]
  PIN timestamp[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 250.280 580.000 250.880 ;
    END
  END timestamp[20]
  PIN timestamp[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 253.000 580.000 253.600 ;
    END
  END timestamp[21]
  PIN timestamp[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 255.720 580.000 256.320 ;
    END
  END timestamp[22]
  PIN timestamp[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 258.440 580.000 259.040 ;
    END
  END timestamp[23]
  PIN timestamp[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 261.160 580.000 261.760 ;
    END
  END timestamp[24]
  PIN timestamp[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 263.880 580.000 264.480 ;
    END
  END timestamp[25]
  PIN timestamp[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 266.600 580.000 267.200 ;
    END
  END timestamp[26]
  PIN timestamp[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 269.320 580.000 269.920 ;
    END
  END timestamp[27]
  PIN timestamp[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 272.040 580.000 272.640 ;
    END
  END timestamp[28]
  PIN timestamp[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 274.760 580.000 275.360 ;
    END
  END timestamp[29]
  PIN timestamp[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 201.320 580.000 201.920 ;
    END
  END timestamp[2]
  PIN timestamp[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 277.480 580.000 278.080 ;
    END
  END timestamp[30]
  PIN timestamp[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 280.200 580.000 280.800 ;
    END
  END timestamp[31]
  PIN timestamp[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 282.920 580.000 283.520 ;
    END
  END timestamp[32]
  PIN timestamp[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 285.640 580.000 286.240 ;
    END
  END timestamp[33]
  PIN timestamp[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 288.360 580.000 288.960 ;
    END
  END timestamp[34]
  PIN timestamp[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 291.080 580.000 291.680 ;
    END
  END timestamp[35]
  PIN timestamp[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 293.800 580.000 294.400 ;
    END
  END timestamp[36]
  PIN timestamp[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 296.520 580.000 297.120 ;
    END
  END timestamp[37]
  PIN timestamp[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 299.240 580.000 299.840 ;
    END
  END timestamp[38]
  PIN timestamp[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 301.960 580.000 302.560 ;
    END
  END timestamp[39]
  PIN timestamp[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 204.040 580.000 204.640 ;
    END
  END timestamp[3]
  PIN timestamp[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 304.680 580.000 305.280 ;
    END
  END timestamp[40]
  PIN timestamp[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 307.400 580.000 308.000 ;
    END
  END timestamp[41]
  PIN timestamp[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 310.120 580.000 310.720 ;
    END
  END timestamp[42]
  PIN timestamp[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 312.840 580.000 313.440 ;
    END
  END timestamp[43]
  PIN timestamp[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 315.560 580.000 316.160 ;
    END
  END timestamp[44]
  PIN timestamp[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 318.280 580.000 318.880 ;
    END
  END timestamp[45]
  PIN timestamp[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 321.000 580.000 321.600 ;
    END
  END timestamp[46]
  PIN timestamp[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 323.720 580.000 324.320 ;
    END
  END timestamp[47]
  PIN timestamp[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 326.440 580.000 327.040 ;
    END
  END timestamp[48]
  PIN timestamp[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 329.160 580.000 329.760 ;
    END
  END timestamp[49]
  PIN timestamp[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 206.760 580.000 207.360 ;
    END
  END timestamp[4]
  PIN timestamp[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 331.880 580.000 332.480 ;
    END
  END timestamp[50]
  PIN timestamp[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 334.600 580.000 335.200 ;
    END
  END timestamp[51]
  PIN timestamp[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 337.320 580.000 337.920 ;
    END
  END timestamp[52]
  PIN timestamp[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 340.040 580.000 340.640 ;
    END
  END timestamp[53]
  PIN timestamp[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 342.760 580.000 343.360 ;
    END
  END timestamp[54]
  PIN timestamp[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 345.480 580.000 346.080 ;
    END
  END timestamp[55]
  PIN timestamp[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 348.200 580.000 348.800 ;
    END
  END timestamp[56]
  PIN timestamp[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 350.920 580.000 351.520 ;
    END
  END timestamp[57]
  PIN timestamp[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 353.640 580.000 354.240 ;
    END
  END timestamp[58]
  PIN timestamp[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 356.360 580.000 356.960 ;
    END
  END timestamp[59]
  PIN timestamp[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 209.480 580.000 210.080 ;
    END
  END timestamp[5]
  PIN timestamp[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 359.080 580.000 359.680 ;
    END
  END timestamp[60]
  PIN timestamp[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 361.800 580.000 362.400 ;
    END
  END timestamp[61]
  PIN timestamp[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 364.520 580.000 365.120 ;
    END
  END timestamp[62]
  PIN timestamp[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 367.240 580.000 367.840 ;
    END
  END timestamp[63]
  PIN timestamp[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 212.200 580.000 212.800 ;
    END
  END timestamp[6]
  PIN timestamp[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 214.920 580.000 215.520 ;
    END
  END timestamp[7]
  PIN timestamp[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 217.640 580.000 218.240 ;
    END
  END timestamp[8]
  PIN timestamp[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 576.000 220.360 580.000 220.960 ;
    END
  END timestamp[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 574.270 568.670 ;
      LAYER li1 ;
        RECT 5.520 10.795 574.080 568.565 ;
      LAYER met1 ;
        RECT 5.520 7.860 575.390 568.720 ;
      LAYER met2 ;
        RECT 7.460 575.720 14.530 576.000 ;
        RECT 15.370 575.720 35.690 576.000 ;
        RECT 36.530 575.720 576.750 576.000 ;
        RECT 7.460 7.830 576.750 575.720 ;
      LAYER met3 ;
        RECT 15.245 498.800 576.775 568.645 ;
        RECT 15.245 497.400 575.600 498.800 ;
        RECT 15.245 496.080 576.775 497.400 ;
        RECT 15.245 494.680 575.600 496.080 ;
        RECT 15.245 493.360 576.775 494.680 ;
        RECT 15.245 491.960 575.600 493.360 ;
        RECT 15.245 490.640 576.775 491.960 ;
        RECT 15.245 489.240 575.600 490.640 ;
        RECT 15.245 487.920 576.775 489.240 ;
        RECT 15.245 486.520 575.600 487.920 ;
        RECT 15.245 485.200 576.775 486.520 ;
        RECT 15.245 483.800 575.600 485.200 ;
        RECT 15.245 482.480 576.775 483.800 ;
        RECT 15.245 481.080 575.600 482.480 ;
        RECT 15.245 479.760 576.775 481.080 ;
        RECT 15.245 478.360 575.600 479.760 ;
        RECT 15.245 477.040 576.775 478.360 ;
        RECT 15.245 475.640 575.600 477.040 ;
        RECT 15.245 474.320 576.775 475.640 ;
        RECT 15.245 472.920 575.600 474.320 ;
        RECT 15.245 471.600 576.775 472.920 ;
        RECT 15.245 470.200 575.600 471.600 ;
        RECT 15.245 468.880 576.775 470.200 ;
        RECT 15.245 467.480 575.600 468.880 ;
        RECT 15.245 466.160 576.775 467.480 ;
        RECT 15.245 464.760 575.600 466.160 ;
        RECT 15.245 463.440 576.775 464.760 ;
        RECT 15.245 462.040 575.600 463.440 ;
        RECT 15.245 460.720 576.775 462.040 ;
        RECT 15.245 459.320 575.600 460.720 ;
        RECT 15.245 458.000 576.775 459.320 ;
        RECT 15.245 456.600 575.600 458.000 ;
        RECT 15.245 455.280 576.775 456.600 ;
        RECT 15.245 453.880 575.600 455.280 ;
        RECT 15.245 452.560 576.775 453.880 ;
        RECT 15.245 451.160 575.600 452.560 ;
        RECT 15.245 449.840 576.775 451.160 ;
        RECT 15.245 448.440 575.600 449.840 ;
        RECT 15.245 447.120 576.775 448.440 ;
        RECT 15.245 445.720 575.600 447.120 ;
        RECT 15.245 444.400 576.775 445.720 ;
        RECT 15.245 443.000 575.600 444.400 ;
        RECT 15.245 441.680 576.775 443.000 ;
        RECT 15.245 440.280 575.600 441.680 ;
        RECT 15.245 438.960 576.775 440.280 ;
        RECT 15.245 437.560 575.600 438.960 ;
        RECT 15.245 436.240 576.775 437.560 ;
        RECT 15.245 434.840 575.600 436.240 ;
        RECT 15.245 433.520 576.775 434.840 ;
        RECT 15.245 432.120 575.600 433.520 ;
        RECT 15.245 430.800 576.775 432.120 ;
        RECT 15.245 429.400 575.600 430.800 ;
        RECT 15.245 428.080 576.775 429.400 ;
        RECT 15.245 426.680 575.600 428.080 ;
        RECT 15.245 425.360 576.775 426.680 ;
        RECT 15.245 423.960 575.600 425.360 ;
        RECT 15.245 422.640 576.775 423.960 ;
        RECT 15.245 421.240 575.600 422.640 ;
        RECT 15.245 419.920 576.775 421.240 ;
        RECT 15.245 418.520 575.600 419.920 ;
        RECT 15.245 417.200 576.775 418.520 ;
        RECT 15.245 415.800 575.600 417.200 ;
        RECT 15.245 414.480 576.775 415.800 ;
        RECT 15.245 413.080 575.600 414.480 ;
        RECT 15.245 411.760 576.775 413.080 ;
        RECT 15.245 410.360 575.600 411.760 ;
        RECT 15.245 409.040 576.775 410.360 ;
        RECT 15.245 407.640 575.600 409.040 ;
        RECT 15.245 406.320 576.775 407.640 ;
        RECT 15.245 404.920 575.600 406.320 ;
        RECT 15.245 403.600 576.775 404.920 ;
        RECT 15.245 402.200 575.600 403.600 ;
        RECT 15.245 400.880 576.775 402.200 ;
        RECT 15.245 399.480 575.600 400.880 ;
        RECT 15.245 398.160 576.775 399.480 ;
        RECT 15.245 396.760 575.600 398.160 ;
        RECT 15.245 395.440 576.775 396.760 ;
        RECT 15.245 394.040 575.600 395.440 ;
        RECT 15.245 392.720 576.775 394.040 ;
        RECT 15.245 391.320 575.600 392.720 ;
        RECT 15.245 390.000 576.775 391.320 ;
        RECT 15.245 388.600 575.600 390.000 ;
        RECT 15.245 387.280 576.775 388.600 ;
        RECT 15.245 385.880 575.600 387.280 ;
        RECT 15.245 384.560 576.775 385.880 ;
        RECT 15.245 383.160 575.600 384.560 ;
        RECT 15.245 381.840 576.775 383.160 ;
        RECT 15.245 380.440 575.600 381.840 ;
        RECT 15.245 379.120 576.775 380.440 ;
        RECT 15.245 377.720 575.600 379.120 ;
        RECT 15.245 376.400 576.775 377.720 ;
        RECT 15.245 375.000 575.600 376.400 ;
        RECT 15.245 373.680 576.775 375.000 ;
        RECT 15.245 372.280 575.600 373.680 ;
        RECT 15.245 370.960 576.775 372.280 ;
        RECT 15.245 369.560 575.600 370.960 ;
        RECT 15.245 368.240 576.775 369.560 ;
        RECT 15.245 366.840 575.600 368.240 ;
        RECT 15.245 365.520 576.775 366.840 ;
        RECT 15.245 364.120 575.600 365.520 ;
        RECT 15.245 362.800 576.775 364.120 ;
        RECT 15.245 361.400 575.600 362.800 ;
        RECT 15.245 360.080 576.775 361.400 ;
        RECT 15.245 358.680 575.600 360.080 ;
        RECT 15.245 357.360 576.775 358.680 ;
        RECT 15.245 355.960 575.600 357.360 ;
        RECT 15.245 354.640 576.775 355.960 ;
        RECT 15.245 353.240 575.600 354.640 ;
        RECT 15.245 351.920 576.775 353.240 ;
        RECT 15.245 350.520 575.600 351.920 ;
        RECT 15.245 349.200 576.775 350.520 ;
        RECT 15.245 347.800 575.600 349.200 ;
        RECT 15.245 346.480 576.775 347.800 ;
        RECT 15.245 345.080 575.600 346.480 ;
        RECT 15.245 343.760 576.775 345.080 ;
        RECT 15.245 342.360 575.600 343.760 ;
        RECT 15.245 341.040 576.775 342.360 ;
        RECT 15.245 339.640 575.600 341.040 ;
        RECT 15.245 338.320 576.775 339.640 ;
        RECT 15.245 336.920 575.600 338.320 ;
        RECT 15.245 335.600 576.775 336.920 ;
        RECT 15.245 334.200 575.600 335.600 ;
        RECT 15.245 332.880 576.775 334.200 ;
        RECT 15.245 331.480 575.600 332.880 ;
        RECT 15.245 330.160 576.775 331.480 ;
        RECT 15.245 328.760 575.600 330.160 ;
        RECT 15.245 327.440 576.775 328.760 ;
        RECT 15.245 326.040 575.600 327.440 ;
        RECT 15.245 324.720 576.775 326.040 ;
        RECT 15.245 323.320 575.600 324.720 ;
        RECT 15.245 322.000 576.775 323.320 ;
        RECT 15.245 320.600 575.600 322.000 ;
        RECT 15.245 319.280 576.775 320.600 ;
        RECT 15.245 317.880 575.600 319.280 ;
        RECT 15.245 316.560 576.775 317.880 ;
        RECT 15.245 315.160 575.600 316.560 ;
        RECT 15.245 313.840 576.775 315.160 ;
        RECT 15.245 312.440 575.600 313.840 ;
        RECT 15.245 311.120 576.775 312.440 ;
        RECT 15.245 309.720 575.600 311.120 ;
        RECT 15.245 308.400 576.775 309.720 ;
        RECT 15.245 307.000 575.600 308.400 ;
        RECT 15.245 305.680 576.775 307.000 ;
        RECT 15.245 304.280 575.600 305.680 ;
        RECT 15.245 302.960 576.775 304.280 ;
        RECT 15.245 301.560 575.600 302.960 ;
        RECT 15.245 300.240 576.775 301.560 ;
        RECT 15.245 298.840 575.600 300.240 ;
        RECT 15.245 297.520 576.775 298.840 ;
        RECT 15.245 296.120 575.600 297.520 ;
        RECT 15.245 294.800 576.775 296.120 ;
        RECT 15.245 293.400 575.600 294.800 ;
        RECT 15.245 292.080 576.775 293.400 ;
        RECT 15.245 290.680 575.600 292.080 ;
        RECT 15.245 289.360 576.775 290.680 ;
        RECT 15.245 287.960 575.600 289.360 ;
        RECT 15.245 286.640 576.775 287.960 ;
        RECT 15.245 285.240 575.600 286.640 ;
        RECT 15.245 283.920 576.775 285.240 ;
        RECT 15.245 282.520 575.600 283.920 ;
        RECT 15.245 281.200 576.775 282.520 ;
        RECT 15.245 279.800 575.600 281.200 ;
        RECT 15.245 278.480 576.775 279.800 ;
        RECT 15.245 277.080 575.600 278.480 ;
        RECT 15.245 275.760 576.775 277.080 ;
        RECT 15.245 274.360 575.600 275.760 ;
        RECT 15.245 273.040 576.775 274.360 ;
        RECT 15.245 271.640 575.600 273.040 ;
        RECT 15.245 270.320 576.775 271.640 ;
        RECT 15.245 268.920 575.600 270.320 ;
        RECT 15.245 267.600 576.775 268.920 ;
        RECT 15.245 266.200 575.600 267.600 ;
        RECT 15.245 264.880 576.775 266.200 ;
        RECT 15.245 263.480 575.600 264.880 ;
        RECT 15.245 262.160 576.775 263.480 ;
        RECT 15.245 260.760 575.600 262.160 ;
        RECT 15.245 259.440 576.775 260.760 ;
        RECT 15.245 258.040 575.600 259.440 ;
        RECT 15.245 256.720 576.775 258.040 ;
        RECT 15.245 255.320 575.600 256.720 ;
        RECT 15.245 254.000 576.775 255.320 ;
        RECT 15.245 252.600 575.600 254.000 ;
        RECT 15.245 251.280 576.775 252.600 ;
        RECT 15.245 249.880 575.600 251.280 ;
        RECT 15.245 248.560 576.775 249.880 ;
        RECT 15.245 247.160 575.600 248.560 ;
        RECT 15.245 245.840 576.775 247.160 ;
        RECT 15.245 244.440 575.600 245.840 ;
        RECT 15.245 243.120 576.775 244.440 ;
        RECT 15.245 241.720 575.600 243.120 ;
        RECT 15.245 240.400 576.775 241.720 ;
        RECT 15.245 239.000 575.600 240.400 ;
        RECT 15.245 237.680 576.775 239.000 ;
        RECT 15.245 236.280 575.600 237.680 ;
        RECT 15.245 234.960 576.775 236.280 ;
        RECT 15.245 233.560 575.600 234.960 ;
        RECT 15.245 232.240 576.775 233.560 ;
        RECT 15.245 230.840 575.600 232.240 ;
        RECT 15.245 229.520 576.775 230.840 ;
        RECT 15.245 228.120 575.600 229.520 ;
        RECT 15.245 226.800 576.775 228.120 ;
        RECT 15.245 225.400 575.600 226.800 ;
        RECT 15.245 224.080 576.775 225.400 ;
        RECT 15.245 222.680 575.600 224.080 ;
        RECT 15.245 221.360 576.775 222.680 ;
        RECT 15.245 219.960 575.600 221.360 ;
        RECT 15.245 218.640 576.775 219.960 ;
        RECT 15.245 217.240 575.600 218.640 ;
        RECT 15.245 215.920 576.775 217.240 ;
        RECT 15.245 214.520 575.600 215.920 ;
        RECT 15.245 213.200 576.775 214.520 ;
        RECT 15.245 211.800 575.600 213.200 ;
        RECT 15.245 210.480 576.775 211.800 ;
        RECT 15.245 209.080 575.600 210.480 ;
        RECT 15.245 207.760 576.775 209.080 ;
        RECT 15.245 206.360 575.600 207.760 ;
        RECT 15.245 205.040 576.775 206.360 ;
        RECT 15.245 203.640 575.600 205.040 ;
        RECT 15.245 202.320 576.775 203.640 ;
        RECT 15.245 200.920 575.600 202.320 ;
        RECT 15.245 199.600 576.775 200.920 ;
        RECT 15.245 198.200 575.600 199.600 ;
        RECT 15.245 196.880 576.775 198.200 ;
        RECT 15.245 195.480 575.600 196.880 ;
        RECT 15.245 194.160 576.775 195.480 ;
        RECT 15.245 192.760 575.600 194.160 ;
        RECT 15.245 191.440 576.775 192.760 ;
        RECT 15.245 190.040 575.600 191.440 ;
        RECT 15.245 188.720 576.775 190.040 ;
        RECT 15.245 187.320 575.600 188.720 ;
        RECT 15.245 186.000 576.775 187.320 ;
        RECT 15.245 184.600 575.600 186.000 ;
        RECT 15.245 183.280 576.775 184.600 ;
        RECT 15.245 181.880 575.600 183.280 ;
        RECT 15.245 180.560 576.775 181.880 ;
        RECT 15.245 179.160 575.600 180.560 ;
        RECT 15.245 177.840 576.775 179.160 ;
        RECT 15.245 176.440 575.600 177.840 ;
        RECT 15.245 175.120 576.775 176.440 ;
        RECT 15.245 173.720 575.600 175.120 ;
        RECT 15.245 172.400 576.775 173.720 ;
        RECT 15.245 171.000 575.600 172.400 ;
        RECT 15.245 169.680 576.775 171.000 ;
        RECT 15.245 168.280 575.600 169.680 ;
        RECT 15.245 166.960 576.775 168.280 ;
        RECT 15.245 165.560 575.600 166.960 ;
        RECT 15.245 164.240 576.775 165.560 ;
        RECT 15.245 162.840 575.600 164.240 ;
        RECT 15.245 161.520 576.775 162.840 ;
        RECT 15.245 160.120 575.600 161.520 ;
        RECT 15.245 158.800 576.775 160.120 ;
        RECT 15.245 157.400 575.600 158.800 ;
        RECT 15.245 156.080 576.775 157.400 ;
        RECT 15.245 154.680 575.600 156.080 ;
        RECT 15.245 153.360 576.775 154.680 ;
        RECT 15.245 151.960 575.600 153.360 ;
        RECT 15.245 150.640 576.775 151.960 ;
        RECT 15.245 149.240 575.600 150.640 ;
        RECT 15.245 147.920 576.775 149.240 ;
        RECT 15.245 146.520 575.600 147.920 ;
        RECT 15.245 145.200 576.775 146.520 ;
        RECT 15.245 143.800 575.600 145.200 ;
        RECT 15.245 142.480 576.775 143.800 ;
        RECT 15.245 141.080 575.600 142.480 ;
        RECT 15.245 139.760 576.775 141.080 ;
        RECT 15.245 138.360 575.600 139.760 ;
        RECT 15.245 137.040 576.775 138.360 ;
        RECT 15.245 135.640 575.600 137.040 ;
        RECT 15.245 134.320 576.775 135.640 ;
        RECT 15.245 132.920 575.600 134.320 ;
        RECT 15.245 131.600 576.775 132.920 ;
        RECT 15.245 130.200 575.600 131.600 ;
        RECT 15.245 128.880 576.775 130.200 ;
        RECT 15.245 127.480 575.600 128.880 ;
        RECT 15.245 126.160 576.775 127.480 ;
        RECT 15.245 124.760 575.600 126.160 ;
        RECT 15.245 123.440 576.775 124.760 ;
        RECT 15.245 122.040 575.600 123.440 ;
        RECT 15.245 120.720 576.775 122.040 ;
        RECT 15.245 119.320 575.600 120.720 ;
        RECT 15.245 118.000 576.775 119.320 ;
        RECT 15.245 116.600 575.600 118.000 ;
        RECT 15.245 115.280 576.775 116.600 ;
        RECT 15.245 113.880 575.600 115.280 ;
        RECT 15.245 112.560 576.775 113.880 ;
        RECT 15.245 111.160 575.600 112.560 ;
        RECT 15.245 109.840 576.775 111.160 ;
        RECT 15.245 108.440 575.600 109.840 ;
        RECT 15.245 107.120 576.775 108.440 ;
        RECT 15.245 105.720 575.600 107.120 ;
        RECT 15.245 104.400 576.775 105.720 ;
        RECT 15.245 103.000 575.600 104.400 ;
        RECT 15.245 101.680 576.775 103.000 ;
        RECT 15.245 100.280 575.600 101.680 ;
        RECT 15.245 98.960 576.775 100.280 ;
        RECT 15.245 97.560 575.600 98.960 ;
        RECT 15.245 96.240 576.775 97.560 ;
        RECT 15.245 94.840 575.600 96.240 ;
        RECT 15.245 93.520 576.775 94.840 ;
        RECT 15.245 92.120 575.600 93.520 ;
        RECT 15.245 90.800 576.775 92.120 ;
        RECT 15.245 89.400 575.600 90.800 ;
        RECT 15.245 88.080 576.775 89.400 ;
        RECT 15.245 86.680 575.600 88.080 ;
        RECT 15.245 85.360 576.775 86.680 ;
        RECT 15.245 83.960 575.600 85.360 ;
        RECT 15.245 82.640 576.775 83.960 ;
        RECT 15.245 81.240 575.600 82.640 ;
        RECT 15.245 10.715 576.775 81.240 ;
      LAYER met4 ;
        RECT 19.615 29.415 20.640 559.465 ;
        RECT 23.040 29.415 23.940 559.465 ;
        RECT 26.340 29.415 100.640 559.465 ;
        RECT 103.040 29.415 103.940 559.465 ;
        RECT 106.340 29.415 180.640 559.465 ;
        RECT 183.040 29.415 183.940 559.465 ;
        RECT 186.340 29.415 260.640 559.465 ;
        RECT 263.040 29.415 263.940 559.465 ;
        RECT 266.340 29.415 340.640 559.465 ;
        RECT 343.040 29.415 343.940 559.465 ;
        RECT 346.340 29.415 420.640 559.465 ;
        RECT 423.040 29.415 423.940 559.465 ;
        RECT 426.340 29.415 500.640 559.465 ;
        RECT 503.040 29.415 503.940 559.465 ;
        RECT 506.340 29.415 571.945 559.465 ;
  END
END ctu_can
END LIBRARY

