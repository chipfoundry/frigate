VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_QSPI_XIP_CTRL_AHBL
  CLASS BLOCK ;
  FOREIGN EF_QSPI_XIP_CTRL_AHBL ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 550.000 ;
  PIN HADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 546.000 41.310 550.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 151.430 546.000 151.710 550.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.470 546.000 162.750 550.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.510 546.000 173.790 550.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 184.550 546.000 184.830 550.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.590 546.000 195.870 550.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.630 546.000 206.910 550.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.670 546.000 217.950 550.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 228.710 546.000 228.990 550.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 239.750 546.000 240.030 550.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 250.790 546.000 251.070 550.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 546.000 52.350 550.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 261.830 546.000 262.110 550.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 272.870 546.000 273.150 550.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.910 546.000 284.190 550.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 294.950 546.000 295.230 550.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 546.000 306.270 550.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 546.000 317.310 550.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 546.000 328.350 550.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 546.000 339.390 550.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 546.000 350.430 550.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 546.000 361.470 550.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 63.110 546.000 63.390 550.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 546.000 372.510 550.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 546.000 383.550 550.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.150 546.000 74.430 550.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 85.190 546.000 85.470 550.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.563400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 96.230 546.000 96.510 550.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 107.270 546.000 107.550 550.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 118.310 546.000 118.590 550.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 129.350 546.000 129.630 550.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 140.390 546.000 140.670 550.000 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 7.910 546.000 8.190 550.000 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 449.510 546.000 449.790 550.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 559.910 546.000 560.190 550.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 570.950 546.000 571.230 550.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 581.990 546.000 582.270 550.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 593.030 546.000 593.310 550.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 604.070 546.000 604.350 550.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 615.110 546.000 615.390 550.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 626.150 546.000 626.430 550.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 637.190 546.000 637.470 550.000 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 648.230 546.000 648.510 550.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 659.270 546.000 659.550 550.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 460.550 546.000 460.830 550.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 670.310 546.000 670.590 550.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 681.350 546.000 681.630 550.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 692.390 546.000 692.670 550.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 703.430 546.000 703.710 550.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 714.470 546.000 714.750 550.000 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 725.510 546.000 725.790 550.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 736.550 546.000 736.830 550.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 747.590 546.000 747.870 550.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 758.630 546.000 758.910 550.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 769.670 546.000 769.950 550.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 471.590 546.000 471.870 550.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 780.710 546.000 780.990 550.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 791.750 546.000 792.030 550.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 482.630 546.000 482.910 550.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 493.670 546.000 493.950 550.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 504.710 546.000 504.990 550.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 515.750 546.000 516.030 550.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 526.790 546.000 527.070 550.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 537.830 546.000 538.110 550.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 548.870 546.000 549.150 550.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 427.430 546.000 427.710 550.000 ;
    END
  END HREADY
  PIN HREADYOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 438.470 546.000 438.750 550.000 ;
    END
  END HREADYOUT
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 18.950 546.000 19.230 550.000 ;
    END
  END HRESETn
  PIN HSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.990 546.000 30.270 550.000 ;
    END
  END HSEL
  PIN HTRANS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 546.000 394.590 550.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 405.350 546.000 405.630 550.000 ;
    END
  END HTRANS[1]
  PIN HWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 546.000 416.670 550.000 ;
    END
  END HWRITE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.340 10.640 105.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.340 10.640 185.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.340 10.640 265.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.340 10.640 345.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 10.640 425.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.340 10.640 505.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 584.340 10.640 585.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.340 10.640 665.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.340 10.640 745.940 538.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.680 794.660 28.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 106.680 794.660 108.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 186.680 794.660 188.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 266.680 794.660 268.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 346.680 794.660 348.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 426.680 794.660 428.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 506.680 794.660 508.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.040 10.640 102.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.040 10.640 182.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.040 10.640 342.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 581.040 10.640 582.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.040 10.640 662.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 538.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 794.660 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 95.080 794.660 96.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 175.080 794.660 176.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 255.080 794.660 256.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 335.080 794.660 336.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 415.080 794.660 416.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 495.080 794.660 496.680 ;
    END
  END VPWR
  PIN ce_n
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END ce_n
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END din[0]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END din[1]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END din[2]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END din[3]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END dout[1]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END dout[2]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END dout[3]
  PIN douten[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END douten[0]
  PIN douten[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END douten[1]
  PIN douten[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END douten[2]
  PIN douten[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END douten[3]
  PIN sck
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END sck
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 794.610 538.645 ;
      LAYER li1 ;
        RECT 5.520 10.795 794.420 538.645 ;
      LAYER met1 ;
        RECT 5.520 10.640 794.420 546.680 ;
      LAYER met2 ;
        RECT 8.470 545.720 18.670 546.710 ;
        RECT 19.510 545.720 29.710 546.710 ;
        RECT 30.550 545.720 40.750 546.710 ;
        RECT 41.590 545.720 51.790 546.710 ;
        RECT 52.630 545.720 62.830 546.710 ;
        RECT 63.670 545.720 73.870 546.710 ;
        RECT 74.710 545.720 84.910 546.710 ;
        RECT 85.750 545.720 95.950 546.710 ;
        RECT 96.790 545.720 106.990 546.710 ;
        RECT 107.830 545.720 118.030 546.710 ;
        RECT 118.870 545.720 129.070 546.710 ;
        RECT 129.910 545.720 140.110 546.710 ;
        RECT 140.950 545.720 151.150 546.710 ;
        RECT 151.990 545.720 162.190 546.710 ;
        RECT 163.030 545.720 173.230 546.710 ;
        RECT 174.070 545.720 184.270 546.710 ;
        RECT 185.110 545.720 195.310 546.710 ;
        RECT 196.150 545.720 206.350 546.710 ;
        RECT 207.190 545.720 217.390 546.710 ;
        RECT 218.230 545.720 228.430 546.710 ;
        RECT 229.270 545.720 239.470 546.710 ;
        RECT 240.310 545.720 250.510 546.710 ;
        RECT 251.350 545.720 261.550 546.710 ;
        RECT 262.390 545.720 272.590 546.710 ;
        RECT 273.430 545.720 283.630 546.710 ;
        RECT 284.470 545.720 294.670 546.710 ;
        RECT 295.510 545.720 305.710 546.710 ;
        RECT 306.550 545.720 316.750 546.710 ;
        RECT 317.590 545.720 327.790 546.710 ;
        RECT 328.630 545.720 338.830 546.710 ;
        RECT 339.670 545.720 349.870 546.710 ;
        RECT 350.710 545.720 360.910 546.710 ;
        RECT 361.750 545.720 371.950 546.710 ;
        RECT 372.790 545.720 382.990 546.710 ;
        RECT 383.830 545.720 394.030 546.710 ;
        RECT 394.870 545.720 405.070 546.710 ;
        RECT 405.910 545.720 416.110 546.710 ;
        RECT 416.950 545.720 427.150 546.710 ;
        RECT 427.990 545.720 438.190 546.710 ;
        RECT 439.030 545.720 449.230 546.710 ;
        RECT 450.070 545.720 460.270 546.710 ;
        RECT 461.110 545.720 471.310 546.710 ;
        RECT 472.150 545.720 482.350 546.710 ;
        RECT 483.190 545.720 493.390 546.710 ;
        RECT 494.230 545.720 504.430 546.710 ;
        RECT 505.270 545.720 515.470 546.710 ;
        RECT 516.310 545.720 526.510 546.710 ;
        RECT 527.350 545.720 537.550 546.710 ;
        RECT 538.390 545.720 548.590 546.710 ;
        RECT 549.430 545.720 559.630 546.710 ;
        RECT 560.470 545.720 570.670 546.710 ;
        RECT 571.510 545.720 581.710 546.710 ;
        RECT 582.550 545.720 592.750 546.710 ;
        RECT 593.590 545.720 603.790 546.710 ;
        RECT 604.630 545.720 614.830 546.710 ;
        RECT 615.670 545.720 625.870 546.710 ;
        RECT 626.710 545.720 636.910 546.710 ;
        RECT 637.750 545.720 647.950 546.710 ;
        RECT 648.790 545.720 658.990 546.710 ;
        RECT 659.830 545.720 670.030 546.710 ;
        RECT 670.870 545.720 681.070 546.710 ;
        RECT 681.910 545.720 692.110 546.710 ;
        RECT 692.950 545.720 703.150 546.710 ;
        RECT 703.990 545.720 714.190 546.710 ;
        RECT 715.030 545.720 725.230 546.710 ;
        RECT 726.070 545.720 736.270 546.710 ;
        RECT 737.110 545.720 747.310 546.710 ;
        RECT 748.150 545.720 758.350 546.710 ;
        RECT 759.190 545.720 769.390 546.710 ;
        RECT 770.230 545.720 780.430 546.710 ;
        RECT 781.270 545.720 791.470 546.710 ;
        RECT 792.310 545.720 792.940 546.710 ;
        RECT 7.980 4.280 792.940 545.720 ;
        RECT 7.980 4.000 28.790 4.280 ;
        RECT 29.630 4.000 85.830 4.280 ;
        RECT 86.670 4.000 142.870 4.280 ;
        RECT 143.710 4.000 199.910 4.280 ;
        RECT 200.750 4.000 256.950 4.280 ;
        RECT 257.790 4.000 313.990 4.280 ;
        RECT 314.830 4.000 371.030 4.280 ;
        RECT 371.870 4.000 428.070 4.280 ;
        RECT 428.910 4.000 485.110 4.280 ;
        RECT 485.950 4.000 542.150 4.280 ;
        RECT 542.990 4.000 599.190 4.280 ;
        RECT 600.030 4.000 656.230 4.280 ;
        RECT 657.070 4.000 713.270 4.280 ;
        RECT 714.110 4.000 770.310 4.280 ;
        RECT 771.150 4.000 792.940 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 788.835 538.725 ;
      LAYER met4 ;
        RECT 96.895 15.815 100.640 533.625 ;
        RECT 103.040 15.815 103.940 533.625 ;
        RECT 106.340 15.815 180.640 533.625 ;
        RECT 183.040 15.815 183.940 533.625 ;
        RECT 186.340 15.815 260.640 533.625 ;
        RECT 263.040 15.815 263.940 533.625 ;
        RECT 266.340 15.815 340.640 533.625 ;
        RECT 343.040 15.815 343.940 533.625 ;
        RECT 346.340 15.815 420.640 533.625 ;
        RECT 423.040 15.815 423.940 533.625 ;
        RECT 426.340 15.815 500.640 533.625 ;
        RECT 503.040 15.815 503.940 533.625 ;
        RECT 506.340 15.815 580.640 533.625 ;
        RECT 583.040 15.815 583.940 533.625 ;
        RECT 586.340 15.815 660.640 533.625 ;
        RECT 663.040 15.815 663.940 533.625 ;
        RECT 666.340 15.815 740.640 533.625 ;
        RECT 743.040 15.815 743.940 533.625 ;
        RECT 746.340 15.815 749.505 533.625 ;
  END
END EF_QSPI_XIP_CTRL_AHBL
END LIBRARY

